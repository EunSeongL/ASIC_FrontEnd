module ctrl (
    
);
    
    
endmodule
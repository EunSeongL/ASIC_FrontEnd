`timescale 1ns/1ps

module twf_02_imag #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output signed [BIT_WIDTH-1:0] twf_out
);

wire signed [BIT_WIDTH-1:0] twf_02_out [0:INDEX_WIDTH-1];

assign twf_out = twf_02_out[index];

assign twf_02_out[0] = 0;
assign twf_02_out[1] = 0;
assign twf_02_out[2] = 0;
assign twf_02_out[3] = 0;
assign twf_02_out[4] = 0;
assign twf_02_out[5] = 0;
assign twf_02_out[6] = 0;
assign twf_02_out[7] = 0;
assign twf_02_out[8] = 0;
assign twf_02_out[9] = 0;
assign twf_02_out[10] = 0;
assign twf_02_out[11] = 0;
assign twf_02_out[12] = 0;
assign twf_02_out[13] = 0;
assign twf_02_out[14] = 0;
assign twf_02_out[15] = 0;
assign twf_02_out[16] = 0;
assign twf_02_out[17] = 0;
assign twf_02_out[18] = 0;
assign twf_02_out[19] = 0;
assign twf_02_out[20] = 0;
assign twf_02_out[21] = 0;
assign twf_02_out[22] = 0;
assign twf_02_out[23] = 0;
assign twf_02_out[24] = 0;
assign twf_02_out[25] = 0;
assign twf_02_out[26] = 0;
assign twf_02_out[27] = 0;
assign twf_02_out[28] = 0;
assign twf_02_out[29] = 0;
assign twf_02_out[30] = 0;
assign twf_02_out[31] = 0;
assign twf_02_out[32] = 0;
assign twf_02_out[33] = 0;
assign twf_02_out[34] = 0;
assign twf_02_out[35] = 0;
assign twf_02_out[36] = 0;
assign twf_02_out[37] = 0;
assign twf_02_out[38] = 0;
assign twf_02_out[39] = 0;
assign twf_02_out[40] = 0;
assign twf_02_out[41] = 0;
assign twf_02_out[42] = 0;
assign twf_02_out[43] = 0;
assign twf_02_out[44] = 0;
assign twf_02_out[45] = 0;
assign twf_02_out[46] = 0;
assign twf_02_out[47] = 0;
assign twf_02_out[48] = 0;
assign twf_02_out[49] = 0;
assign twf_02_out[50] = 0;
assign twf_02_out[51] = 0;
assign twf_02_out[52] = 0;
assign twf_02_out[53] = 0;
assign twf_02_out[54] = 0;
assign twf_02_out[55] = 0;
assign twf_02_out[56] = 0;
assign twf_02_out[57] = 0;
assign twf_02_out[58] = 0;
assign twf_02_out[59] = 0;
assign twf_02_out[60] = 0;
assign twf_02_out[61] = 0;
assign twf_02_out[62] = 0;
assign twf_02_out[63] = 0;
assign twf_02_out[64] = 0;
assign twf_02_out[65] = -6;
assign twf_02_out[66] = -13;
assign twf_02_out[67] = -19;
assign twf_02_out[68] = -25;
assign twf_02_out[69] = -31;
assign twf_02_out[70] = -37;
assign twf_02_out[71] = -43;
assign twf_02_out[72] = -49;
assign twf_02_out[73] = -55;
assign twf_02_out[74] = -60;
assign twf_02_out[75] = -66;
assign twf_02_out[76] = -71;
assign twf_02_out[77] = -76;
assign twf_02_out[78] = -81;
assign twf_02_out[79] = -86;
assign twf_02_out[80] = -91;
assign twf_02_out[81] = -95;
assign twf_02_out[82] = -99;
assign twf_02_out[83] = -103;
assign twf_02_out[84] = -106;
assign twf_02_out[85] = -110;
assign twf_02_out[86] = -113;
assign twf_02_out[87] = -116;
assign twf_02_out[88] = -118;
assign twf_02_out[89] = -121;
assign twf_02_out[90] = -122;
assign twf_02_out[91] = -124;
assign twf_02_out[92] = -126;
assign twf_02_out[93] = -127;
assign twf_02_out[94] = -127;
assign twf_02_out[95] = -128;
assign twf_02_out[96] = -128;
assign twf_02_out[97] = -128;
assign twf_02_out[98] = -127;
assign twf_02_out[99] = -127;
assign twf_02_out[100] = -126;
assign twf_02_out[101] = -124;
assign twf_02_out[102] = -122;
assign twf_02_out[103] = -121;
assign twf_02_out[104] = -118;
assign twf_02_out[105] = -116;
assign twf_02_out[106] = -113;
assign twf_02_out[107] = -110;
assign twf_02_out[108] = -106;
assign twf_02_out[109] = -103;
assign twf_02_out[110] = -99;
assign twf_02_out[111] = -95;
assign twf_02_out[112] = -91;
assign twf_02_out[113] = -86;
assign twf_02_out[114] = -81;
assign twf_02_out[115] = -76;
assign twf_02_out[116] = -71;
assign twf_02_out[117] = -66;
assign twf_02_out[118] = -60;
assign twf_02_out[119] = -55;
assign twf_02_out[120] = -49;
assign twf_02_out[121] = -43;
assign twf_02_out[122] = -37;
assign twf_02_out[123] = -31;
assign twf_02_out[124] = -25;
assign twf_02_out[125] = -19;
assign twf_02_out[126] = -13;
assign twf_02_out[127] = -6;
assign twf_02_out[128] = 0;
assign twf_02_out[129] = -3;
assign twf_02_out[130] = -6;
assign twf_02_out[131] = -9;
assign twf_02_out[132] = -13;
assign twf_02_out[133] = -16;
assign twf_02_out[134] = -19;
assign twf_02_out[135] = -22;
assign twf_02_out[136] = -25;
assign twf_02_out[137] = -28;
assign twf_02_out[138] = -31;
assign twf_02_out[139] = -34;
assign twf_02_out[140] = -37;
assign twf_02_out[141] = -40;
assign twf_02_out[142] = -43;
assign twf_02_out[143] = -46;
assign twf_02_out[144] = -49;
assign twf_02_out[145] = -52;
assign twf_02_out[146] = -55;
assign twf_02_out[147] = -58;
assign twf_02_out[148] = -60;
assign twf_02_out[149] = -63;
assign twf_02_out[150] = -66;
assign twf_02_out[151] = -68;
assign twf_02_out[152] = -71;
assign twf_02_out[153] = -74;
assign twf_02_out[154] = -76;
assign twf_02_out[155] = -79;
assign twf_02_out[156] = -81;
assign twf_02_out[157] = -84;
assign twf_02_out[158] = -86;
assign twf_02_out[159] = -88;
assign twf_02_out[160] = -91;
assign twf_02_out[161] = -93;
assign twf_02_out[162] = -95;
assign twf_02_out[163] = -97;
assign twf_02_out[164] = -99;
assign twf_02_out[165] = -101;
assign twf_02_out[166] = -103;
assign twf_02_out[167] = -105;
assign twf_02_out[168] = -106;
assign twf_02_out[169] = -108;
assign twf_02_out[170] = -110;
assign twf_02_out[171] = -111;
assign twf_02_out[172] = -113;
assign twf_02_out[173] = -114;
assign twf_02_out[174] = -116;
assign twf_02_out[175] = -117;
assign twf_02_out[176] = -118;
assign twf_02_out[177] = -119;
assign twf_02_out[178] = -121;
assign twf_02_out[179] = -122;
assign twf_02_out[180] = -122;
assign twf_02_out[181] = -123;
assign twf_02_out[182] = -124;
assign twf_02_out[183] = -125;
assign twf_02_out[184] = -126;
assign twf_02_out[185] = -126;
assign twf_02_out[186] = -127;
assign twf_02_out[187] = -127;
assign twf_02_out[188] = -127;
assign twf_02_out[189] = -128;
assign twf_02_out[190] = -128;
assign twf_02_out[191] = -128;
assign twf_02_out[192] = 0;
assign twf_02_out[193] = -9;
assign twf_02_out[194] = -19;
assign twf_02_out[195] = -28;
assign twf_02_out[196] = -37;
assign twf_02_out[197] = -46;
assign twf_02_out[198] = -55;
assign twf_02_out[199] = -63;
assign twf_02_out[200] = -71;
assign twf_02_out[201] = -79;
assign twf_02_out[202] = -86;
assign twf_02_out[203] = -93;
assign twf_02_out[204] = -99;
assign twf_02_out[205] = -105;
assign twf_02_out[206] = -110;
assign twf_02_out[207] = -114;
assign twf_02_out[208] = -118;
assign twf_02_out[209] = -122;
assign twf_02_out[210] = -124;
assign twf_02_out[211] = -126;
assign twf_02_out[212] = -127;
assign twf_02_out[213] = -128;
assign twf_02_out[214] = -128;
assign twf_02_out[215] = -127;
assign twf_02_out[216] = -126;
assign twf_02_out[217] = -123;
assign twf_02_out[218] = -121;
assign twf_02_out[219] = -117;
assign twf_02_out[220] = -113;
assign twf_02_out[221] = -108;
assign twf_02_out[222] = -103;
assign twf_02_out[223] = -97;
assign twf_02_out[224] = -91;
assign twf_02_out[225] = -84;
assign twf_02_out[226] = -76;
assign twf_02_out[227] = -68;
assign twf_02_out[228] = -60;
assign twf_02_out[229] = -52;
assign twf_02_out[230] = -43;
assign twf_02_out[231] = -34;
assign twf_02_out[232] = -25;
assign twf_02_out[233] = -16;
assign twf_02_out[234] = -6;
assign twf_02_out[235] = 3;
assign twf_02_out[236] = 13;
assign twf_02_out[237] = 22;
assign twf_02_out[238] = 31;
assign twf_02_out[239] = 40;
assign twf_02_out[240] = 49;
assign twf_02_out[241] = 58;
assign twf_02_out[242] = 66;
assign twf_02_out[243] = 74;
assign twf_02_out[244] = 81;
assign twf_02_out[245] = 88;
assign twf_02_out[246] = 95;
assign twf_02_out[247] = 101;
assign twf_02_out[248] = 106;
assign twf_02_out[249] = 111;
assign twf_02_out[250] = 116;
assign twf_02_out[251] = 119;
assign twf_02_out[252] = 122;
assign twf_02_out[253] = 125;
assign twf_02_out[254] = 127;
assign twf_02_out[255] = 128;
assign twf_02_out[256] = 0;
assign twf_02_out[257] = -2;
assign twf_02_out[258] = -3;
assign twf_02_out[259] = -5;
assign twf_02_out[260] = -6;
assign twf_02_out[261] = -8;
assign twf_02_out[262] = -9;
assign twf_02_out[263] = -11;
assign twf_02_out[264] = -13;
assign twf_02_out[265] = -14;
assign twf_02_out[266] = -16;
assign twf_02_out[267] = -17;
assign twf_02_out[268] = -19;
assign twf_02_out[269] = -20;
assign twf_02_out[270] = -22;
assign twf_02_out[271] = -23;
assign twf_02_out[272] = -25;
assign twf_02_out[273] = -27;
assign twf_02_out[274] = -28;
assign twf_02_out[275] = -30;
assign twf_02_out[276] = -31;
assign twf_02_out[277] = -33;
assign twf_02_out[278] = -34;
assign twf_02_out[279] = -36;
assign twf_02_out[280] = -37;
assign twf_02_out[281] = -39;
assign twf_02_out[282] = -40;
assign twf_02_out[283] = -42;
assign twf_02_out[284] = -43;
assign twf_02_out[285] = -45;
assign twf_02_out[286] = -46;
assign twf_02_out[287] = -48;
assign twf_02_out[288] = -49;
assign twf_02_out[289] = -50;
assign twf_02_out[290] = -52;
assign twf_02_out[291] = -53;
assign twf_02_out[292] = -55;
assign twf_02_out[293] = -56;
assign twf_02_out[294] = -58;
assign twf_02_out[295] = -59;
assign twf_02_out[296] = -60;
assign twf_02_out[297] = -62;
assign twf_02_out[298] = -63;
assign twf_02_out[299] = -64;
assign twf_02_out[300] = -66;
assign twf_02_out[301] = -67;
assign twf_02_out[302] = -68;
assign twf_02_out[303] = -70;
assign twf_02_out[304] = -71;
assign twf_02_out[305] = -72;
assign twf_02_out[306] = -74;
assign twf_02_out[307] = -75;
assign twf_02_out[308] = -76;
assign twf_02_out[309] = -78;
assign twf_02_out[310] = -79;
assign twf_02_out[311] = -80;
assign twf_02_out[312] = -81;
assign twf_02_out[313] = -82;
assign twf_02_out[314] = -84;
assign twf_02_out[315] = -85;
assign twf_02_out[316] = -86;
assign twf_02_out[317] = -87;
assign twf_02_out[318] = -88;
assign twf_02_out[319] = -89;
assign twf_02_out[320] = 0;
assign twf_02_out[321] = -8;
assign twf_02_out[322] = -16;
assign twf_02_out[323] = -23;
assign twf_02_out[324] = -31;
assign twf_02_out[325] = -39;
assign twf_02_out[326] = -46;
assign twf_02_out[327] = -53;
assign twf_02_out[328] = -60;
assign twf_02_out[329] = -67;
assign twf_02_out[330] = -74;
assign twf_02_out[331] = -80;
assign twf_02_out[332] = -86;
assign twf_02_out[333] = -92;
assign twf_02_out[334] = -97;
assign twf_02_out[335] = -102;
assign twf_02_out[336] = -106;
assign twf_02_out[337] = -111;
assign twf_02_out[338] = -114;
assign twf_02_out[339] = -118;
assign twf_02_out[340] = -121;
assign twf_02_out[341] = -123;
assign twf_02_out[342] = -125;
assign twf_02_out[343] = -126;
assign twf_02_out[344] = -127;
assign twf_02_out[345] = -128;
assign twf_02_out[346] = -128;
assign twf_02_out[347] = -128;
assign twf_02_out[348] = -127;
assign twf_02_out[349] = -125;
assign twf_02_out[350] = -123;
assign twf_02_out[351] = -121;
assign twf_02_out[352] = -118;
assign twf_02_out[353] = -115;
assign twf_02_out[354] = -111;
assign twf_02_out[355] = -107;
assign twf_02_out[356] = -103;
assign twf_02_out[357] = -98;
assign twf_02_out[358] = -93;
assign twf_02_out[359] = -87;
assign twf_02_out[360] = -81;
assign twf_02_out[361] = -75;
assign twf_02_out[362] = -68;
assign twf_02_out[363] = -62;
assign twf_02_out[364] = -55;
assign twf_02_out[365] = -48;
assign twf_02_out[366] = -40;
assign twf_02_out[367] = -33;
assign twf_02_out[368] = -25;
assign twf_02_out[369] = -17;
assign twf_02_out[370] = -9;
assign twf_02_out[371] = -2;
assign twf_02_out[372] = 6;
assign twf_02_out[373] = 14;
assign twf_02_out[374] = 22;
assign twf_02_out[375] = 30;
assign twf_02_out[376] = 37;
assign twf_02_out[377] = 45;
assign twf_02_out[378] = 52;
assign twf_02_out[379] = 59;
assign twf_02_out[380] = 66;
assign twf_02_out[381] = 72;
assign twf_02_out[382] = 79;
assign twf_02_out[383] = 85;
assign twf_02_out[384] = 0;
assign twf_02_out[385] = -5;
assign twf_02_out[386] = -9;
assign twf_02_out[387] = -14;
assign twf_02_out[388] = -19;
assign twf_02_out[389] = -23;
assign twf_02_out[390] = -28;
assign twf_02_out[391] = -33;
assign twf_02_out[392] = -37;
assign twf_02_out[393] = -42;
assign twf_02_out[394] = -46;
assign twf_02_out[395] = -50;
assign twf_02_out[396] = -55;
assign twf_02_out[397] = -59;
assign twf_02_out[398] = -63;
assign twf_02_out[399] = -67;
assign twf_02_out[400] = -71;
assign twf_02_out[401] = -75;
assign twf_02_out[402] = -79;
assign twf_02_out[403] = -82;
assign twf_02_out[404] = -86;
assign twf_02_out[405] = -89;
assign twf_02_out[406] = -93;
assign twf_02_out[407] = -96;
assign twf_02_out[408] = -99;
assign twf_02_out[409] = -102;
assign twf_02_out[410] = -105;
assign twf_02_out[411] = -107;
assign twf_02_out[412] = -110;
assign twf_02_out[413] = -112;
assign twf_02_out[414] = -114;
assign twf_02_out[415] = -116;
assign twf_02_out[416] = -118;
assign twf_02_out[417] = -120;
assign twf_02_out[418] = -122;
assign twf_02_out[419] = -123;
assign twf_02_out[420] = -124;
assign twf_02_out[421] = -125;
assign twf_02_out[422] = -126;
assign twf_02_out[423] = -127;
assign twf_02_out[424] = -127;
assign twf_02_out[425] = -128;
assign twf_02_out[426] = -128;
assign twf_02_out[427] = -128;
assign twf_02_out[428] = -128;
assign twf_02_out[429] = -128;
assign twf_02_out[430] = -127;
assign twf_02_out[431] = -126;
assign twf_02_out[432] = -126;
assign twf_02_out[433] = -125;
assign twf_02_out[434] = -123;
assign twf_02_out[435] = -122;
assign twf_02_out[436] = -121;
assign twf_02_out[437] = -119;
assign twf_02_out[438] = -117;
assign twf_02_out[439] = -115;
assign twf_02_out[440] = -113;
assign twf_02_out[441] = -111;
assign twf_02_out[442] = -108;
assign twf_02_out[443] = -106;
assign twf_02_out[444] = -103;
assign twf_02_out[445] = -100;
assign twf_02_out[446] = -97;
assign twf_02_out[447] = -94;
assign twf_02_out[448] = 0;
assign twf_02_out[449] = -11;
assign twf_02_out[450] = -22;
assign twf_02_out[451] = -33;
assign twf_02_out[452] = -43;
assign twf_02_out[453] = -53;
assign twf_02_out[454] = -63;
assign twf_02_out[455] = -72;
assign twf_02_out[456] = -81;
assign twf_02_out[457] = -89;
assign twf_02_out[458] = -97;
assign twf_02_out[459] = -104;
assign twf_02_out[460] = -110;
assign twf_02_out[461] = -115;
assign twf_02_out[462] = -119;
assign twf_02_out[463] = -123;
assign twf_02_out[464] = -126;
assign twf_02_out[465] = -127;
assign twf_02_out[466] = -128;
assign twf_02_out[467] = -128;
assign twf_02_out[468] = -127;
assign twf_02_out[469] = -125;
assign twf_02_out[470] = -122;
assign twf_02_out[471] = -118;
assign twf_02_out[472] = -113;
assign twf_02_out[473] = -107;
assign twf_02_out[474] = -101;
assign twf_02_out[475] = -94;
assign twf_02_out[476] = -86;
assign twf_02_out[477] = -78;
assign twf_02_out[478] = -68;
assign twf_02_out[479] = -59;
assign twf_02_out[480] = -49;
assign twf_02_out[481] = -39;
assign twf_02_out[482] = -28;
assign twf_02_out[483] = -17;
assign twf_02_out[484] = -6;
assign twf_02_out[485] = 5;
assign twf_02_out[486] = 16;
assign twf_02_out[487] = 27;
assign twf_02_out[488] = 37;
assign twf_02_out[489] = 48;
assign twf_02_out[490] = 58;
assign twf_02_out[491] = 67;
assign twf_02_out[492] = 76;
assign twf_02_out[493] = 85;
assign twf_02_out[494] = 93;
assign twf_02_out[495] = 100;
assign twf_02_out[496] = 106;
assign twf_02_out[497] = 112;
assign twf_02_out[498] = 117;
assign twf_02_out[499] = 121;
assign twf_02_out[500] = 124;
assign twf_02_out[501] = 126;
assign twf_02_out[502] = 128;
assign twf_02_out[503] = 128;
assign twf_02_out[504] = 127;
assign twf_02_out[505] = 126;
assign twf_02_out[506] = 123;
assign twf_02_out[507] = 120;
assign twf_02_out[508] = 116;
assign twf_02_out[509] = 111;
assign twf_02_out[510] = 105;
assign twf_02_out[511] = 98;

endmodule

`timescale 1ns/1ps

module twf_02_imag #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output logic signed [BIT_WIDTH-1:0] twf_out
);

always @(*) begin
    case(index)
        0: twf_out = 0;
        1: twf_out = 0;
        2: twf_out = 0;
        3: twf_out = 0;
        4: twf_out = 0;
        5: twf_out = 0;
        6: twf_out = 0;
        7: twf_out = 0;
        8: twf_out = 0;
        9: twf_out = 0;
        10: twf_out = 0;
        11: twf_out = 0;
        12: twf_out = 0;
        13: twf_out = 0;
        14: twf_out = 0;
        15: twf_out = 0;
        16: twf_out = 0;
        17: twf_out = 0;
        18: twf_out = 0;
        19: twf_out = 0;
        20: twf_out = 0;
        21: twf_out = 0;
        22: twf_out = 0;
        23: twf_out = 0;
        24: twf_out = 0;
        25: twf_out = 0;
        26: twf_out = 0;
        27: twf_out = 0;
        28: twf_out = 0;
        29: twf_out = 0;
        30: twf_out = 0;
        31: twf_out = 0;
        32: twf_out = 0;
        33: twf_out = 0;
        34: twf_out = 0;
        35: twf_out = 0;
        36: twf_out = 0;
        37: twf_out = 0;
        38: twf_out = 0;
        39: twf_out = 0;
        40: twf_out = 0;
        41: twf_out = 0;
        42: twf_out = 0;
        43: twf_out = 0;
        44: twf_out = 0;
        45: twf_out = 0;
        46: twf_out = 0;
        47: twf_out = 0;
        48: twf_out = 0;
        49: twf_out = 0;
        50: twf_out = 0;
        51: twf_out = 0;
        52: twf_out = 0;
        53: twf_out = 0;
        54: twf_out = 0;
        55: twf_out = 0;
        56: twf_out = 0;
        57: twf_out = 0;
        58: twf_out = 0;
        59: twf_out = 0;
        60: twf_out = 0;
        61: twf_out = 0;
        62: twf_out = 0;
        63: twf_out = 0;
        64: twf_out = 0;
        65: twf_out = -6;
        66: twf_out = -13;
        67: twf_out = -19;
        68: twf_out = -25;
        69: twf_out = -31;
        70: twf_out = -37;
        71: twf_out = -43;
        72: twf_out = -49;
        73: twf_out = -55;
        74: twf_out = -60;
        75: twf_out = -66;
        76: twf_out = -71;
        77: twf_out = -76;
        78: twf_out = -81;
        79: twf_out = -86;
        80: twf_out = -91;
        81: twf_out = -95;
        82: twf_out = -99;
        83: twf_out = -103;
        84: twf_out = -106;
        85: twf_out = -110;
        86: twf_out = -113;
        87: twf_out = -116;
        88: twf_out = -118;
        89: twf_out = -121;
        90: twf_out = -122;
        91: twf_out = -124;
        92: twf_out = -126;
        93: twf_out = -127;
        94: twf_out = -127;
        95: twf_out = -128;
        96: twf_out = -128;
        97: twf_out = -128;
        98: twf_out = -127;
        99: twf_out = -127;
        100: twf_out = -126;
        101: twf_out = -124;
        102: twf_out = -122;
        103: twf_out = -121;
        104: twf_out = -118;
        105: twf_out = -116;
        106: twf_out = -113;
        107: twf_out = -110;
        108: twf_out = -106;
        109: twf_out = -103;
        110: twf_out = -99;
        111: twf_out = -95;
        112: twf_out = -91;
        113: twf_out = -86;
        114: twf_out = -81;
        115: twf_out = -76;
        116: twf_out = -71;
        117: twf_out = -66;
        118: twf_out = -60;
        119: twf_out = -55;
        120: twf_out = -49;
        121: twf_out = -43;
        122: twf_out = -37;
        123: twf_out = -31;
        124: twf_out = -25;
        125: twf_out = -19;
        126: twf_out = -13;
        127: twf_out = -6;
        128: twf_out = 0;
        129: twf_out = -3;
        130: twf_out = -6;
        131: twf_out = -9;
        132: twf_out = -13;
        133: twf_out = -16;
        134: twf_out = -19;
        135: twf_out = -22;
        136: twf_out = -25;
        137: twf_out = -28;
        138: twf_out = -31;
        139: twf_out = -34;
        140: twf_out = -37;
        141: twf_out = -40;
        142: twf_out = -43;
        143: twf_out = -46;
        144: twf_out = -49;
        145: twf_out = -52;
        146: twf_out = -55;
        147: twf_out = -58;
        148: twf_out = -60;
        149: twf_out = -63;
        150: twf_out = -66;
        151: twf_out = -68;
        152: twf_out = -71;
        153: twf_out = -74;
        154: twf_out = -76;
        155: twf_out = -79;
        156: twf_out = -81;
        157: twf_out = -84;
        158: twf_out = -86;
        159: twf_out = -88;
        160: twf_out = -91;
        161: twf_out = -93;
        162: twf_out = -95;
        163: twf_out = -97;
        164: twf_out = -99;
        165: twf_out = -101;
        166: twf_out = -103;
        167: twf_out = -105;
        168: twf_out = -106;
        169: twf_out = -108;
        170: twf_out = -110;
        171: twf_out = -111;
        172: twf_out = -113;
        173: twf_out = -114;
        174: twf_out = -116;
        175: twf_out = -117;
        176: twf_out = -118;
        177: twf_out = -119;
        178: twf_out = -121;
        179: twf_out = -122;
        180: twf_out = -122;
        181: twf_out = -123;
        182: twf_out = -124;
        183: twf_out = -125;
        184: twf_out = -126;
        185: twf_out = -126;
        186: twf_out = -127;
        187: twf_out = -127;
        188: twf_out = -127;
        189: twf_out = -128;
        190: twf_out = -128;
        191: twf_out = -128;
        192: twf_out = 0;
        193: twf_out = -9;
        194: twf_out = -19;
        195: twf_out = -28;
        196: twf_out = -37;
        197: twf_out = -46;
        198: twf_out = -55;
        199: twf_out = -63;
        200: twf_out = -71;
        201: twf_out = -79;
        202: twf_out = -86;
        203: twf_out = -93;
        204: twf_out = -99;
        205: twf_out = -105;
        206: twf_out = -110;
        207: twf_out = -114;
        208: twf_out = -118;
        209: twf_out = -122;
        210: twf_out = -124;
        211: twf_out = -126;
        212: twf_out = -127;
        213: twf_out = -128;
        214: twf_out = -128;
        215: twf_out = -127;
        216: twf_out = -126;
        217: twf_out = -123;
        218: twf_out = -121;
        219: twf_out = -117;
        220: twf_out = -113;
        221: twf_out = -108;
        222: twf_out = -103;
        223: twf_out = -97;
        224: twf_out = -91;
        225: twf_out = -84;
        226: twf_out = -76;
        227: twf_out = -68;
        228: twf_out = -60;
        229: twf_out = -52;
        230: twf_out = -43;
        231: twf_out = -34;
        232: twf_out = -25;
        233: twf_out = -16;
        234: twf_out = -6;
        235: twf_out = 3;
        236: twf_out = 13;
        237: twf_out = 22;
        238: twf_out = 31;
        239: twf_out = 40;
        240: twf_out = 49;
        241: twf_out = 58;
        242: twf_out = 66;
        243: twf_out = 74;
        244: twf_out = 81;
        245: twf_out = 88;
        246: twf_out = 95;
        247: twf_out = 101;
        248: twf_out = 106;
        249: twf_out = 111;
        250: twf_out = 116;
        251: twf_out = 119;
        252: twf_out = 122;
        253: twf_out = 125;
        254: twf_out = 127;
        255: twf_out = 128;
        256: twf_out = 0;
        257: twf_out = -2;
        258: twf_out = -3;
        259: twf_out = -5;
        260: twf_out = -6;
        261: twf_out = -8;
        262: twf_out = -9;
        263: twf_out = -11;
        264: twf_out = -13;
        265: twf_out = -14;
        266: twf_out = -16;
        267: twf_out = -17;
        268: twf_out = -19;
        269: twf_out = -20;
        270: twf_out = -22;
        271: twf_out = -23;
        272: twf_out = -25;
        273: twf_out = -27;
        274: twf_out = -28;
        275: twf_out = -30;
        276: twf_out = -31;
        277: twf_out = -33;
        278: twf_out = -34;
        279: twf_out = -36;
        280: twf_out = -37;
        281: twf_out = -39;
        282: twf_out = -40;
        283: twf_out = -42;
        284: twf_out = -43;
        285: twf_out = -45;
        286: twf_out = -46;
        287: twf_out = -48;
        288: twf_out = -49;
        289: twf_out = -50;
        290: twf_out = -52;
        291: twf_out = -53;
        292: twf_out = -55;
        293: twf_out = -56;
        294: twf_out = -58;
        295: twf_out = -59;
        296: twf_out = -60;
        297: twf_out = -62;
        298: twf_out = -63;
        299: twf_out = -64;
        300: twf_out = -66;
        301: twf_out = -67;
        302: twf_out = -68;
        303: twf_out = -70;
        304: twf_out = -71;
        305: twf_out = -72;
        306: twf_out = -74;
        307: twf_out = -75;
        308: twf_out = -76;
        309: twf_out = -78;
        310: twf_out = -79;
        311: twf_out = -80;
        312: twf_out = -81;
        313: twf_out = -82;
        314: twf_out = -84;
        315: twf_out = -85;
        316: twf_out = -86;
        317: twf_out = -87;
        318: twf_out = -88;
        319: twf_out = -89;
        320: twf_out = 0;
        321: twf_out = -8;
        322: twf_out = -16;
        323: twf_out = -23;
        324: twf_out = -31;
        325: twf_out = -39;
        326: twf_out = -46;
        327: twf_out = -53;
        328: twf_out = -60;
        329: twf_out = -67;
        330: twf_out = -74;
        331: twf_out = -80;
        332: twf_out = -86;
        333: twf_out = -92;
        334: twf_out = -97;
        335: twf_out = -102;
        336: twf_out = -106;
        337: twf_out = -111;
        338: twf_out = -114;
        339: twf_out = -118;
        340: twf_out = -121;
        341: twf_out = -123;
        342: twf_out = -125;
        343: twf_out = -126;
        344: twf_out = -127;
        345: twf_out = -128;
        346: twf_out = -128;
        347: twf_out = -128;
        348: twf_out = -127;
        349: twf_out = -125;
        350: twf_out = -123;
        351: twf_out = -121;
        352: twf_out = -118;
        353: twf_out = -115;
        354: twf_out = -111;
        355: twf_out = -107;
        356: twf_out = -103;
        357: twf_out = -98;
        358: twf_out = -93;
        359: twf_out = -87;
        360: twf_out = -81;
        361: twf_out = -75;
        362: twf_out = -68;
        363: twf_out = -62;
        364: twf_out = -55;
        365: twf_out = -48;
        366: twf_out = -40;
        367: twf_out = -33;
        368: twf_out = -25;
        369: twf_out = -17;
        370: twf_out = -9;
        371: twf_out = -2;
        372: twf_out = 6;
        373: twf_out = 14;
        374: twf_out = 22;
        375: twf_out = 30;
        376: twf_out = 37;
        377: twf_out = 45;
        378: twf_out = 52;
        379: twf_out = 59;
        380: twf_out = 66;
        381: twf_out = 72;
        382: twf_out = 79;
        383: twf_out = 85;
        384: twf_out = 0;
        385: twf_out = -5;
        386: twf_out = -9;
        387: twf_out = -14;
        388: twf_out = -19;
        389: twf_out = -23;
        390: twf_out = -28;
        391: twf_out = -33;
        392: twf_out = -37;
        393: twf_out = -42;
        394: twf_out = -46;
        395: twf_out = -50;
        396: twf_out = -55;
        397: twf_out = -59;
        398: twf_out = -63;
        399: twf_out = -67;
        400: twf_out = -71;
        401: twf_out = -75;
        402: twf_out = -79;
        403: twf_out = -82;
        404: twf_out = -86;
        405: twf_out = -89;
        406: twf_out = -93;
        407: twf_out = -96;
        408: twf_out = -99;
        409: twf_out = -102;
        410: twf_out = -105;
        411: twf_out = -107;
        412: twf_out = -110;
        413: twf_out = -112;
        414: twf_out = -114;
        415: twf_out = -116;
        416: twf_out = -118;
        417: twf_out = -120;
        418: twf_out = -122;
        419: twf_out = -123;
        420: twf_out = -124;
        421: twf_out = -125;
        422: twf_out = -126;
        423: twf_out = -127;
        424: twf_out = -127;
        425: twf_out = -128;
        426: twf_out = -128;
        427: twf_out = -128;
        428: twf_out = -128;
        429: twf_out = -128;
        430: twf_out = -127;
        431: twf_out = -126;
        432: twf_out = -126;
        433: twf_out = -125;
        434: twf_out = -123;
        435: twf_out = -122;
        436: twf_out = -121;
        437: twf_out = -119;
        438: twf_out = -117;
        439: twf_out = -115;
        440: twf_out = -113;
        441: twf_out = -111;
        442: twf_out = -108;
        443: twf_out = -106;
        444: twf_out = -103;
        445: twf_out = -100;
        446: twf_out = -97;
        447: twf_out = -94;
        448: twf_out = 0;
        449: twf_out = -11;
        450: twf_out = -22;
        451: twf_out = -33;
        452: twf_out = -43;
        453: twf_out = -53;
        454: twf_out = -63;
        455: twf_out = -72;
        456: twf_out = -81;
        457: twf_out = -89;
        458: twf_out = -97;
        459: twf_out = -104;
        460: twf_out = -110;
        461: twf_out = -115;
        462: twf_out = -119;
        463: twf_out = -123;
        464: twf_out = -126;
        465: twf_out = -127;
        466: twf_out = -128;
        467: twf_out = -128;
        468: twf_out = -127;
        469: twf_out = -125;
        470: twf_out = -122;
        471: twf_out = -118;
        472: twf_out = -113;
        473: twf_out = -107;
        474: twf_out = -101;
        475: twf_out = -94;
        476: twf_out = -86;
        477: twf_out = -78;
        478: twf_out = -68;
        479: twf_out = -59;
        480: twf_out = -49;
        481: twf_out = -39;
        482: twf_out = -28;
        483: twf_out = -17;
        484: twf_out = -6;
        485: twf_out = 5;
        486: twf_out = 16;
        487: twf_out = 27;
        488: twf_out = 37;
        489: twf_out = 48;
        490: twf_out = 58;
        491: twf_out = 67;
        492: twf_out = 76;
        493: twf_out = 85;
        494: twf_out = 93;
        495: twf_out = 100;
        496: twf_out = 106;
        497: twf_out = 112;
        498: twf_out = 117;
        499: twf_out = 121;
        500: twf_out = 124;
        501: twf_out = 126;
        502: twf_out = 128;
        503: twf_out = 128;
        504: twf_out = 127;
        505: twf_out = 126;
        506: twf_out = 123;
        507: twf_out = 120;
        508: twf_out = 116;
        509: twf_out = 111;
        510: twf_out = 105;
        511: twf_out = 98;
        default: twf_out = 0;
    endcase
end

endmodule

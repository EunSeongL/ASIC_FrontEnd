`timescale 1ns/1ps

module step02_twf #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output logic signed [BIT_WIDTH-1:0] twf_out
);

always @(*) begin
    case(index)
        0: twf_out = 128;
        1: twf_out = 128;
        2: twf_out = 128;
        3: twf_out = 128;
        4: twf_out = 128;
        5: twf_out = 128;
        6: twf_out = 128;
        7: twf_out = 128;
        8: twf_out = 128;
        9: twf_out = 128;
        10: twf_out = 128;
        11: twf_out = 128;
        12: twf_out = 128;
        13: twf_out = 128;
        14: twf_out = 128;
        15: twf_out = 128;
        16: twf_out = 128;
        17: twf_out = 128;
        18: twf_out = 128;
        19: twf_out = 128;
        20: twf_out = 128;
        21: twf_out = 128;
        22: twf_out = 128;
        23: twf_out = 128;
        24: twf_out = 128;
        25: twf_out = 128;
        26: twf_out = 128;
        27: twf_out = 128;
        28: twf_out = 128;
        29: twf_out = 128;
        30: twf_out = 128;
        31: twf_out = 128;
        32: twf_out = 128;
        33: twf_out = 128;
        34: twf_out = 128;
        35: twf_out = 128;
        36: twf_out = 128;
        37: twf_out = 128;
        38: twf_out = 128;
        39: twf_out = 128;
        40: twf_out = 128;
        41: twf_out = 128;
        42: twf_out = 128;
        43: twf_out = 128;
        44: twf_out = 128;
        45: twf_out = 128;
        46: twf_out = 128;
        47: twf_out = 128;
        48: twf_out = 128;
        49: twf_out = 128;
        50: twf_out = 128;
        51: twf_out = 128;
        52: twf_out = 128;
        53: twf_out = 128;
        54: twf_out = 128;
        55: twf_out = 128;
        56: twf_out = 128;
        57: twf_out = 128;
        58: twf_out = 128;
        59: twf_out = 128;
        60: twf_out = 128;
        61: twf_out = 128;
        62: twf_out = 128;
        63: twf_out = 128;
        64: twf_out = 128;
        65: twf_out = 128;
        66: twf_out = 127;
        67: twf_out = 127;
        68: twf_out = 126;
        69: twf_out = 124;
        70: twf_out = 122;
        71: twf_out = 121;
        72: twf_out = 118;
        73: twf_out = 116;
        74: twf_out = 113;
        75: twf_out = 110;
        76: twf_out = 106;
        77: twf_out = 103;
        78: twf_out = 99;
        79: twf_out = 95;
        80: twf_out = 91;
        81: twf_out = 86;
        82: twf_out = 81;
        83: twf_out = 76;
        84: twf_out = 71;
        85: twf_out = 66;
        86: twf_out = 60;
        87: twf_out = 55;
        88: twf_out = 49;
        89: twf_out = 43;
        90: twf_out = 37;
        91: twf_out = 31;
        92: twf_out = 25;
        93: twf_out = 19;
        94: twf_out = 13;
        95: twf_out = 6;
        96: twf_out = 0;
        97: twf_out = -6;
        98: twf_out = -13;
        99: twf_out = -19;
        100: twf_out = -25;
        101: twf_out = -31;
        102: twf_out = -37;
        103: twf_out = -43;
        104: twf_out = -49;
        105: twf_out = -55;
        106: twf_out = -60;
        107: twf_out = -66;
        108: twf_out = -71;
        109: twf_out = -76;
        110: twf_out = -81;
        111: twf_out = -86;
        112: twf_out = -91;
        113: twf_out = -95;
        114: twf_out = -99;
        115: twf_out = -103;
        116: twf_out = -106;
        117: twf_out = -110;
        118: twf_out = -113;
        119: twf_out = -116;
        120: twf_out = -118;
        121: twf_out = -121;
        122: twf_out = -122;
        123: twf_out = -124;
        124: twf_out = -126;
        125: twf_out = -127;
        126: twf_out = -127;
        127: twf_out = -128;
        128: twf_out = 128;
        129: twf_out = 128;
        130: twf_out = 128;
        131: twf_out = 128;
        132: twf_out = 127;
        133: twf_out = 127;
        134: twf_out = 127;
        135: twf_out = 126;
        136: twf_out = 126;
        137: twf_out = 125;
        138: twf_out = 124;
        139: twf_out = 123;
        140: twf_out = 122;
        141: twf_out = 122;
        142: twf_out = 121;
        143: twf_out = 119;
        144: twf_out = 118;
        145: twf_out = 117;
        146: twf_out = 116;
        147: twf_out = 114;
        148: twf_out = 113;
        149: twf_out = 111;
        150: twf_out = 110;
        151: twf_out = 108;
        152: twf_out = 106;
        153: twf_out = 105;
        154: twf_out = 103;
        155: twf_out = 101;
        156: twf_out = 99;
        157: twf_out = 97;
        158: twf_out = 95;
        159: twf_out = 93;
        160: twf_out = 91;
        161: twf_out = 88;
        162: twf_out = 86;
        163: twf_out = 84;
        164: twf_out = 81;
        165: twf_out = 79;
        166: twf_out = 76;
        167: twf_out = 74;
        168: twf_out = 71;
        169: twf_out = 68;
        170: twf_out = 66;
        171: twf_out = 63;
        172: twf_out = 60;
        173: twf_out = 58;
        174: twf_out = 55;
        175: twf_out = 52;
        176: twf_out = 49;
        177: twf_out = 46;
        178: twf_out = 43;
        179: twf_out = 40;
        180: twf_out = 37;
        181: twf_out = 34;
        182: twf_out = 31;
        183: twf_out = 28;
        184: twf_out = 25;
        185: twf_out = 22;
        186: twf_out = 19;
        187: twf_out = 16;
        188: twf_out = 13;
        189: twf_out = 9;
        190: twf_out = 6;
        191: twf_out = 3;
        192: twf_out = 128;
        193: twf_out = 128;
        194: twf_out = 127;
        195: twf_out = 125;
        196: twf_out = 122;
        197: twf_out = 119;
        198: twf_out = 116;
        199: twf_out = 111;
        200: twf_out = 106;
        201: twf_out = 101;
        202: twf_out = 95;
        203: twf_out = 88;
        204: twf_out = 81;
        205: twf_out = 74;
        206: twf_out = 66;
        207: twf_out = 58;
        208: twf_out = 49;
        209: twf_out = 40;
        210: twf_out = 31;
        211: twf_out = 22;
        212: twf_out = 13;
        213: twf_out = 3;
        214: twf_out = -6;
        215: twf_out = -16;
        216: twf_out = -25;
        217: twf_out = -34;
        218: twf_out = -43;
        219: twf_out = -52;
        220: twf_out = -60;
        221: twf_out = -68;
        222: twf_out = -76;
        223: twf_out = -84;
        224: twf_out = -91;
        225: twf_out = -97;
        226: twf_out = -103;
        227: twf_out = -108;
        228: twf_out = -113;
        229: twf_out = -117;
        230: twf_out = -121;
        231: twf_out = -123;
        232: twf_out = -126;
        233: twf_out = -127;
        234: twf_out = -128;
        235: twf_out = -128;
        236: twf_out = -127;
        237: twf_out = -126;
        238: twf_out = -124;
        239: twf_out = -122;
        240: twf_out = -118;
        241: twf_out = -114;
        242: twf_out = -110;
        243: twf_out = -105;
        244: twf_out = -99;
        245: twf_out = -93;
        246: twf_out = -86;
        247: twf_out = -79;
        248: twf_out = -71;
        249: twf_out = -63;
        250: twf_out = -55;
        251: twf_out = -46;
        252: twf_out = -37;
        253: twf_out = -28;
        254: twf_out = -19;
        255: twf_out = -9;
        256: twf_out = 128;
        257: twf_out = 128;
        258: twf_out = 128;
        259: twf_out = 128;
        260: twf_out = 128;
        261: twf_out = 128;
        262: twf_out = 128;
        263: twf_out = 128;
        264: twf_out = 127;
        265: twf_out = 127;
        266: twf_out = 127;
        267: twf_out = 127;
        268: twf_out = 127;
        269: twf_out = 126;
        270: twf_out = 126;
        271: twf_out = 126;
        272: twf_out = 126;
        273: twf_out = 125;
        274: twf_out = 125;
        275: twf_out = 125;
        276: twf_out = 124;
        277: twf_out = 124;
        278: twf_out = 123;
        279: twf_out = 123;
        280: twf_out = 122;
        281: twf_out = 122;
        282: twf_out = 122;
        283: twf_out = 121;
        284: twf_out = 121;
        285: twf_out = 120;
        286: twf_out = 119;
        287: twf_out = 119;
        288: twf_out = 118;
        289: twf_out = 118;
        290: twf_out = 117;
        291: twf_out = 116;
        292: twf_out = 116;
        293: twf_out = 115;
        294: twf_out = 114;
        295: twf_out = 114;
        296: twf_out = 113;
        297: twf_out = 112;
        298: twf_out = 111;
        299: twf_out = 111;
        300: twf_out = 110;
        301: twf_out = 109;
        302: twf_out = 108;
        303: twf_out = 107;
        304: twf_out = 106;
        305: twf_out = 106;
        306: twf_out = 105;
        307: twf_out = 104;
        308: twf_out = 103;
        309: twf_out = 102;
        310: twf_out = 101;
        311: twf_out = 100;
        312: twf_out = 99;
        313: twf_out = 98;
        314: twf_out = 97;
        315: twf_out = 96;
        316: twf_out = 95;
        317: twf_out = 94;
        318: twf_out = 93;
        319: twf_out = 92;
        320: twf_out = 128;
        321: twf_out = 128;
        322: twf_out = 127;
        323: twf_out = 126;
        324: twf_out = 124;
        325: twf_out = 122;
        326: twf_out = 119;
        327: twf_out = 116;
        328: twf_out = 113;
        329: twf_out = 109;
        330: twf_out = 105;
        331: twf_out = 100;
        332: twf_out = 95;
        333: twf_out = 89;
        334: twf_out = 84;
        335: twf_out = 78;
        336: twf_out = 71;
        337: twf_out = 64;
        338: twf_out = 58;
        339: twf_out = 50;
        340: twf_out = 43;
        341: twf_out = 36;
        342: twf_out = 28;
        343: twf_out = 20;
        344: twf_out = 13;
        345: twf_out = 5;
        346: twf_out = -3;
        347: twf_out = -11;
        348: twf_out = -19;
        349: twf_out = -27;
        350: twf_out = -34;
        351: twf_out = -42;
        352: twf_out = -49;
        353: twf_out = -56;
        354: twf_out = -63;
        355: twf_out = -70;
        356: twf_out = -76;
        357: twf_out = -82;
        358: twf_out = -88;
        359: twf_out = -94;
        360: twf_out = -99;
        361: twf_out = -104;
        362: twf_out = -108;
        363: twf_out = -112;
        364: twf_out = -116;
        365: twf_out = -119;
        366: twf_out = -122;
        367: twf_out = -124;
        368: twf_out = -126;
        369: twf_out = -127;
        370: twf_out = -128;
        371: twf_out = -128;
        372: twf_out = -128;
        373: twf_out = -127;
        374: twf_out = -126;
        375: twf_out = -125;
        376: twf_out = -122;
        377: twf_out = -120;
        378: twf_out = -117;
        379: twf_out = -114;
        380: twf_out = -110;
        381: twf_out = -106;
        382: twf_out = -101;
        383: twf_out = -96;
        384: twf_out = 128;
        385: twf_out = 128;
        386: twf_out = 128;
        387: twf_out = 127;
        388: twf_out = 127;
        389: twf_out = 126;
        390: twf_out = 125;
        391: twf_out = 124;
        392: twf_out = 122;
        393: twf_out = 121;
        394: twf_out = 119;
        395: twf_out = 118;
        396: twf_out = 116;
        397: twf_out = 114;
        398: twf_out = 111;
        399: twf_out = 109;
        400: twf_out = 106;
        401: twf_out = 104;
        402: twf_out = 101;
        403: twf_out = 98;
        404: twf_out = 95;
        405: twf_out = 92;
        406: twf_out = 88;
        407: twf_out = 85;
        408: twf_out = 81;
        409: twf_out = 78;
        410: twf_out = 74;
        411: twf_out = 70;
        412: twf_out = 66;
        413: twf_out = 62;
        414: twf_out = 58;
        415: twf_out = 53;
        416: twf_out = 49;
        417: twf_out = 45;
        418: twf_out = 40;
        419: twf_out = 36;
        420: twf_out = 31;
        421: twf_out = 27;
        422: twf_out = 22;
        423: twf_out = 17;
        424: twf_out = 13;
        425: twf_out = 8;
        426: twf_out = 3;
        427: twf_out = -2;
        428: twf_out = -6;
        429: twf_out = -11;
        430: twf_out = -16;
        431: twf_out = -20;
        432: twf_out = -25;
        433: twf_out = -30;
        434: twf_out = -34;
        435: twf_out = -39;
        436: twf_out = -43;
        437: twf_out = -48;
        438: twf_out = -52;
        439: twf_out = -56;
        440: twf_out = -60;
        441: twf_out = -64;
        442: twf_out = -68;
        443: twf_out = -72;
        444: twf_out = -76;
        445: twf_out = -80;
        446: twf_out = -84;
        447: twf_out = -87;
        448: twf_out = 128;
        449: twf_out = 128;
        450: twf_out = 126;
        451: twf_out = 124;
        452: twf_out = 121;
        453: twf_out = 116;
        454: twf_out = 111;
        455: twf_out = 106;
        456: twf_out = 99;
        457: twf_out = 92;
        458: twf_out = 84;
        459: twf_out = 75;
        460: twf_out = 66;
        461: twf_out = 56;
        462: twf_out = 46;
        463: twf_out = 36;
        464: twf_out = 25;
        465: twf_out = 14;
        466: twf_out = 3;
        467: twf_out = -8;
        468: twf_out = -19;
        469: twf_out = -30;
        470: twf_out = -40;
        471: twf_out = -50;
        472: twf_out = -60;
        473: twf_out = -70;
        474: twf_out = -79;
        475: twf_out = -87;
        476: twf_out = -95;
        477: twf_out = -102;
        478: twf_out = -108;
        479: twf_out = -114;
        480: twf_out = -118;
        481: twf_out = -122;
        482: twf_out = -125;
        483: twf_out = -127;
        484: twf_out = -128;
        485: twf_out = -128;
        486: twf_out = -127;
        487: twf_out = -125;
        488: twf_out = -122;
        489: twf_out = -119;
        490: twf_out = -114;
        491: twf_out = -109;
        492: twf_out = -103;
        493: twf_out = -96;
        494: twf_out = -88;
        495: twf_out = -80;
        496: twf_out = -71;
        497: twf_out = -62;
        498: twf_out = -52;
        499: twf_out = -42;
        500: twf_out = -31;
        501: twf_out = -20;
        502: twf_out = -9;
        503: twf_out = 2;
        504: twf_out = 13;
        505: twf_out = 23;
        506: twf_out = 34;
        507: twf_out = 45;
        508: twf_out = 55;
        509: twf_out = 64;
        510: twf_out = 74;
        511: twf_out = 82;
        default: twf_out = 0;
    endcase
end

endmodule

`timescale 1ns/1ps

module twf_12_real #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output signed [BIT_WIDTH-1:0] twf_out
);

wire signed [BIT_WIDTH-1:0] twf_12_out [0:INDEX_WIDTH-1];

assign twf_out = twf_12_out[index];

assign twf_12_out[0] = 128;
assign twf_12_out[1] = 128;
assign twf_12_out[2] = 128;
assign twf_12_out[3] = 128;
assign twf_12_out[4] = 128;
assign twf_12_out[5] = 128;
assign twf_12_out[6] = 128;
assign twf_12_out[7] = 128;
assign twf_12_out[8] = 128;
assign twf_12_out[9] = 118;
assign twf_12_out[10] = 91;
assign twf_12_out[11] = 49;
assign twf_12_out[12] = 0;
assign twf_12_out[13] = -49;
assign twf_12_out[14] = -91;
assign twf_12_out[15] = -118;
assign twf_12_out[16] = 128;
assign twf_12_out[17] = 126;
assign twf_12_out[18] = 118;
assign twf_12_out[19] = 106;
assign twf_12_out[20] = 91;
assign twf_12_out[21] = 71;
assign twf_12_out[22] = 49;
assign twf_12_out[23] = 25;
assign twf_12_out[24] = 128;
assign twf_12_out[25] = 106;
assign twf_12_out[26] = 49;
assign twf_12_out[27] = -25;
assign twf_12_out[28] = -91;
assign twf_12_out[29] = -126;
assign twf_12_out[30] = -118;
assign twf_12_out[31] = -71;
assign twf_12_out[32] = 128;
assign twf_12_out[33] = 127;
assign twf_12_out[34] = 126;
assign twf_12_out[35] = 122;
assign twf_12_out[36] = 118;
assign twf_12_out[37] = 113;
assign twf_12_out[38] = 106;
assign twf_12_out[39] = 99;
assign twf_12_out[40] = 128;
assign twf_12_out[41] = 113;
assign twf_12_out[42] = 71;
assign twf_12_out[43] = 13;
assign twf_12_out[44] = -49;
assign twf_12_out[45] = -99;
assign twf_12_out[46] = -126;
assign twf_12_out[47] = -122;
assign twf_12_out[48] = 128;
assign twf_12_out[49] = 122;
assign twf_12_out[50] = 106;
assign twf_12_out[51] = 81;
assign twf_12_out[52] = 49;
assign twf_12_out[53] = 13;
assign twf_12_out[54] = -25;
assign twf_12_out[55] = -60;
assign twf_12_out[56] = 128;
assign twf_12_out[57] = 99;
assign twf_12_out[58] = 25;
assign twf_12_out[59] = -60;
assign twf_12_out[60] = -118;
assign twf_12_out[61] = -122;
assign twf_12_out[62] = -71;
assign twf_12_out[63] = 13;
assign twf_12_out[64] = 128;
assign twf_12_out[65] = 128;
assign twf_12_out[66] = 128;
assign twf_12_out[67] = 128;
assign twf_12_out[68] = 128;
assign twf_12_out[69] = 128;
assign twf_12_out[70] = 128;
assign twf_12_out[71] = 128;
assign twf_12_out[72] = 128;
assign twf_12_out[73] = 118;
assign twf_12_out[74] = 91;
assign twf_12_out[75] = 49;
assign twf_12_out[76] = 0;
assign twf_12_out[77] = -49;
assign twf_12_out[78] = -91;
assign twf_12_out[79] = -118;
assign twf_12_out[80] = 128;
assign twf_12_out[81] = 126;
assign twf_12_out[82] = 118;
assign twf_12_out[83] = 106;
assign twf_12_out[84] = 91;
assign twf_12_out[85] = 71;
assign twf_12_out[86] = 49;
assign twf_12_out[87] = 25;
assign twf_12_out[88] = 128;
assign twf_12_out[89] = 106;
assign twf_12_out[90] = 49;
assign twf_12_out[91] = -25;
assign twf_12_out[92] = -91;
assign twf_12_out[93] = -126;
assign twf_12_out[94] = -118;
assign twf_12_out[95] = -71;
assign twf_12_out[96] = 128;
assign twf_12_out[97] = 127;
assign twf_12_out[98] = 126;
assign twf_12_out[99] = 122;
assign twf_12_out[100] = 118;
assign twf_12_out[101] = 113;
assign twf_12_out[102] = 106;
assign twf_12_out[103] = 99;
assign twf_12_out[104] = 128;
assign twf_12_out[105] = 113;
assign twf_12_out[106] = 71;
assign twf_12_out[107] = 13;
assign twf_12_out[108] = -49;
assign twf_12_out[109] = -99;
assign twf_12_out[110] = -126;
assign twf_12_out[111] = -122;
assign twf_12_out[112] = 128;
assign twf_12_out[113] = 122;
assign twf_12_out[114] = 106;
assign twf_12_out[115] = 81;
assign twf_12_out[116] = 49;
assign twf_12_out[117] = 13;
assign twf_12_out[118] = -25;
assign twf_12_out[119] = -60;
assign twf_12_out[120] = 128;
assign twf_12_out[121] = 99;
assign twf_12_out[122] = 25;
assign twf_12_out[123] = -60;
assign twf_12_out[124] = -118;
assign twf_12_out[125] = -122;
assign twf_12_out[126] = -71;
assign twf_12_out[127] = 13;
assign twf_12_out[128] = 128;
assign twf_12_out[129] = 128;
assign twf_12_out[130] = 128;
assign twf_12_out[131] = 128;
assign twf_12_out[132] = 128;
assign twf_12_out[133] = 128;
assign twf_12_out[134] = 128;
assign twf_12_out[135] = 128;
assign twf_12_out[136] = 128;
assign twf_12_out[137] = 118;
assign twf_12_out[138] = 91;
assign twf_12_out[139] = 49;
assign twf_12_out[140] = 0;
assign twf_12_out[141] = -49;
assign twf_12_out[142] = -91;
assign twf_12_out[143] = -118;
assign twf_12_out[144] = 128;
assign twf_12_out[145] = 126;
assign twf_12_out[146] = 118;
assign twf_12_out[147] = 106;
assign twf_12_out[148] = 91;
assign twf_12_out[149] = 71;
assign twf_12_out[150] = 49;
assign twf_12_out[151] = 25;
assign twf_12_out[152] = 128;
assign twf_12_out[153] = 106;
assign twf_12_out[154] = 49;
assign twf_12_out[155] = -25;
assign twf_12_out[156] = -91;
assign twf_12_out[157] = -126;
assign twf_12_out[158] = -118;
assign twf_12_out[159] = -71;
assign twf_12_out[160] = 128;
assign twf_12_out[161] = 127;
assign twf_12_out[162] = 126;
assign twf_12_out[163] = 122;
assign twf_12_out[164] = 118;
assign twf_12_out[165] = 113;
assign twf_12_out[166] = 106;
assign twf_12_out[167] = 99;
assign twf_12_out[168] = 128;
assign twf_12_out[169] = 113;
assign twf_12_out[170] = 71;
assign twf_12_out[171] = 13;
assign twf_12_out[172] = -49;
assign twf_12_out[173] = -99;
assign twf_12_out[174] = -126;
assign twf_12_out[175] = -122;
assign twf_12_out[176] = 128;
assign twf_12_out[177] = 122;
assign twf_12_out[178] = 106;
assign twf_12_out[179] = 81;
assign twf_12_out[180] = 49;
assign twf_12_out[181] = 13;
assign twf_12_out[182] = -25;
assign twf_12_out[183] = -60;
assign twf_12_out[184] = 128;
assign twf_12_out[185] = 99;
assign twf_12_out[186] = 25;
assign twf_12_out[187] = -60;
assign twf_12_out[188] = -118;
assign twf_12_out[189] = -122;
assign twf_12_out[190] = -71;
assign twf_12_out[191] = 13;
assign twf_12_out[192] = 128;
assign twf_12_out[193] = 128;
assign twf_12_out[194] = 128;
assign twf_12_out[195] = 128;
assign twf_12_out[196] = 128;
assign twf_12_out[197] = 128;
assign twf_12_out[198] = 128;
assign twf_12_out[199] = 128;
assign twf_12_out[200] = 128;
assign twf_12_out[201] = 118;
assign twf_12_out[202] = 91;
assign twf_12_out[203] = 49;
assign twf_12_out[204] = 0;
assign twf_12_out[205] = -49;
assign twf_12_out[206] = -91;
assign twf_12_out[207] = -118;
assign twf_12_out[208] = 128;
assign twf_12_out[209] = 126;
assign twf_12_out[210] = 118;
assign twf_12_out[211] = 106;
assign twf_12_out[212] = 91;
assign twf_12_out[213] = 71;
assign twf_12_out[214] = 49;
assign twf_12_out[215] = 25;
assign twf_12_out[216] = 128;
assign twf_12_out[217] = 106;
assign twf_12_out[218] = 49;
assign twf_12_out[219] = -25;
assign twf_12_out[220] = -91;
assign twf_12_out[221] = -126;
assign twf_12_out[222] = -118;
assign twf_12_out[223] = -71;
assign twf_12_out[224] = 128;
assign twf_12_out[225] = 127;
assign twf_12_out[226] = 126;
assign twf_12_out[227] = 122;
assign twf_12_out[228] = 118;
assign twf_12_out[229] = 113;
assign twf_12_out[230] = 106;
assign twf_12_out[231] = 99;
assign twf_12_out[232] = 128;
assign twf_12_out[233] = 113;
assign twf_12_out[234] = 71;
assign twf_12_out[235] = 13;
assign twf_12_out[236] = -49;
assign twf_12_out[237] = -99;
assign twf_12_out[238] = -126;
assign twf_12_out[239] = -122;
assign twf_12_out[240] = 128;
assign twf_12_out[241] = 122;
assign twf_12_out[242] = 106;
assign twf_12_out[243] = 81;
assign twf_12_out[244] = 49;
assign twf_12_out[245] = 13;
assign twf_12_out[246] = -25;
assign twf_12_out[247] = -60;
assign twf_12_out[248] = 128;
assign twf_12_out[249] = 99;
assign twf_12_out[250] = 25;
assign twf_12_out[251] = -60;
assign twf_12_out[252] = -118;
assign twf_12_out[253] = -122;
assign twf_12_out[254] = -71;
assign twf_12_out[255] = 13;
assign twf_12_out[256] = 128;
assign twf_12_out[257] = 128;
assign twf_12_out[258] = 128;
assign twf_12_out[259] = 128;
assign twf_12_out[260] = 128;
assign twf_12_out[261] = 128;
assign twf_12_out[262] = 128;
assign twf_12_out[263] = 128;
assign twf_12_out[264] = 128;
assign twf_12_out[265] = 118;
assign twf_12_out[266] = 91;
assign twf_12_out[267] = 49;
assign twf_12_out[268] = 0;
assign twf_12_out[269] = -49;
assign twf_12_out[270] = -91;
assign twf_12_out[271] = -118;
assign twf_12_out[272] = 128;
assign twf_12_out[273] = 126;
assign twf_12_out[274] = 118;
assign twf_12_out[275] = 106;
assign twf_12_out[276] = 91;
assign twf_12_out[277] = 71;
assign twf_12_out[278] = 49;
assign twf_12_out[279] = 25;
assign twf_12_out[280] = 128;
assign twf_12_out[281] = 106;
assign twf_12_out[282] = 49;
assign twf_12_out[283] = -25;
assign twf_12_out[284] = -91;
assign twf_12_out[285] = -126;
assign twf_12_out[286] = -118;
assign twf_12_out[287] = -71;
assign twf_12_out[288] = 128;
assign twf_12_out[289] = 127;
assign twf_12_out[290] = 126;
assign twf_12_out[291] = 122;
assign twf_12_out[292] = 118;
assign twf_12_out[293] = 113;
assign twf_12_out[294] = 106;
assign twf_12_out[295] = 99;
assign twf_12_out[296] = 128;
assign twf_12_out[297] = 113;
assign twf_12_out[298] = 71;
assign twf_12_out[299] = 13;
assign twf_12_out[300] = -49;
assign twf_12_out[301] = -99;
assign twf_12_out[302] = -126;
assign twf_12_out[303] = -122;
assign twf_12_out[304] = 128;
assign twf_12_out[305] = 122;
assign twf_12_out[306] = 106;
assign twf_12_out[307] = 81;
assign twf_12_out[308] = 49;
assign twf_12_out[309] = 13;
assign twf_12_out[310] = -25;
assign twf_12_out[311] = -60;
assign twf_12_out[312] = 128;
assign twf_12_out[313] = 99;
assign twf_12_out[314] = 25;
assign twf_12_out[315] = -60;
assign twf_12_out[316] = -118;
assign twf_12_out[317] = -122;
assign twf_12_out[318] = -71;
assign twf_12_out[319] = 13;
assign twf_12_out[320] = 128;
assign twf_12_out[321] = 128;
assign twf_12_out[322] = 128;
assign twf_12_out[323] = 128;
assign twf_12_out[324] = 128;
assign twf_12_out[325] = 128;
assign twf_12_out[326] = 128;
assign twf_12_out[327] = 128;
assign twf_12_out[328] = 128;
assign twf_12_out[329] = 118;
assign twf_12_out[330] = 91;
assign twf_12_out[331] = 49;
assign twf_12_out[332] = 0;
assign twf_12_out[333] = -49;
assign twf_12_out[334] = -91;
assign twf_12_out[335] = -118;
assign twf_12_out[336] = 128;
assign twf_12_out[337] = 126;
assign twf_12_out[338] = 118;
assign twf_12_out[339] = 106;
assign twf_12_out[340] = 91;
assign twf_12_out[341] = 71;
assign twf_12_out[342] = 49;
assign twf_12_out[343] = 25;
assign twf_12_out[344] = 128;
assign twf_12_out[345] = 106;
assign twf_12_out[346] = 49;
assign twf_12_out[347] = -25;
assign twf_12_out[348] = -91;
assign twf_12_out[349] = -126;
assign twf_12_out[350] = -118;
assign twf_12_out[351] = -71;
assign twf_12_out[352] = 128;
assign twf_12_out[353] = 127;
assign twf_12_out[354] = 126;
assign twf_12_out[355] = 122;
assign twf_12_out[356] = 118;
assign twf_12_out[357] = 113;
assign twf_12_out[358] = 106;
assign twf_12_out[359] = 99;
assign twf_12_out[360] = 128;
assign twf_12_out[361] = 113;
assign twf_12_out[362] = 71;
assign twf_12_out[363] = 13;
assign twf_12_out[364] = -49;
assign twf_12_out[365] = -99;
assign twf_12_out[366] = -126;
assign twf_12_out[367] = -122;
assign twf_12_out[368] = 128;
assign twf_12_out[369] = 122;
assign twf_12_out[370] = 106;
assign twf_12_out[371] = 81;
assign twf_12_out[372] = 49;
assign twf_12_out[373] = 13;
assign twf_12_out[374] = -25;
assign twf_12_out[375] = -60;
assign twf_12_out[376] = 128;
assign twf_12_out[377] = 99;
assign twf_12_out[378] = 25;
assign twf_12_out[379] = -60;
assign twf_12_out[380] = -118;
assign twf_12_out[381] = -122;
assign twf_12_out[382] = -71;
assign twf_12_out[383] = 13;
assign twf_12_out[384] = 128;
assign twf_12_out[385] = 128;
assign twf_12_out[386] = 128;
assign twf_12_out[387] = 128;
assign twf_12_out[388] = 128;
assign twf_12_out[389] = 128;
assign twf_12_out[390] = 128;
assign twf_12_out[391] = 128;
assign twf_12_out[392] = 128;
assign twf_12_out[393] = 118;
assign twf_12_out[394] = 91;
assign twf_12_out[395] = 49;
assign twf_12_out[396] = 0;
assign twf_12_out[397] = -49;
assign twf_12_out[398] = -91;
assign twf_12_out[399] = -118;
assign twf_12_out[400] = 128;
assign twf_12_out[401] = 126;
assign twf_12_out[402] = 118;
assign twf_12_out[403] = 106;
assign twf_12_out[404] = 91;
assign twf_12_out[405] = 71;
assign twf_12_out[406] = 49;
assign twf_12_out[407] = 25;
assign twf_12_out[408] = 128;
assign twf_12_out[409] = 106;
assign twf_12_out[410] = 49;
assign twf_12_out[411] = -25;
assign twf_12_out[412] = -91;
assign twf_12_out[413] = -126;
assign twf_12_out[414] = -118;
assign twf_12_out[415] = -71;
assign twf_12_out[416] = 128;
assign twf_12_out[417] = 127;
assign twf_12_out[418] = 126;
assign twf_12_out[419] = 122;
assign twf_12_out[420] = 118;
assign twf_12_out[421] = 113;
assign twf_12_out[422] = 106;
assign twf_12_out[423] = 99;
assign twf_12_out[424] = 128;
assign twf_12_out[425] = 113;
assign twf_12_out[426] = 71;
assign twf_12_out[427] = 13;
assign twf_12_out[428] = -49;
assign twf_12_out[429] = -99;
assign twf_12_out[430] = -126;
assign twf_12_out[431] = -122;
assign twf_12_out[432] = 128;
assign twf_12_out[433] = 122;
assign twf_12_out[434] = 106;
assign twf_12_out[435] = 81;
assign twf_12_out[436] = 49;
assign twf_12_out[437] = 13;
assign twf_12_out[438] = -25;
assign twf_12_out[439] = -60;
assign twf_12_out[440] = 128;
assign twf_12_out[441] = 99;
assign twf_12_out[442] = 25;
assign twf_12_out[443] = -60;
assign twf_12_out[444] = -118;
assign twf_12_out[445] = -122;
assign twf_12_out[446] = -71;
assign twf_12_out[447] = 13;
assign twf_12_out[448] = 128;
assign twf_12_out[449] = 128;
assign twf_12_out[450] = 128;
assign twf_12_out[451] = 128;
assign twf_12_out[452] = 128;
assign twf_12_out[453] = 128;
assign twf_12_out[454] = 128;
assign twf_12_out[455] = 128;
assign twf_12_out[456] = 128;
assign twf_12_out[457] = 118;
assign twf_12_out[458] = 91;
assign twf_12_out[459] = 49;
assign twf_12_out[460] = 0;
assign twf_12_out[461] = -49;
assign twf_12_out[462] = -91;
assign twf_12_out[463] = -118;
assign twf_12_out[464] = 128;
assign twf_12_out[465] = 126;
assign twf_12_out[466] = 118;
assign twf_12_out[467] = 106;
assign twf_12_out[468] = 91;
assign twf_12_out[469] = 71;
assign twf_12_out[470] = 49;
assign twf_12_out[471] = 25;
assign twf_12_out[472] = 128;
assign twf_12_out[473] = 106;
assign twf_12_out[474] = 49;
assign twf_12_out[475] = -25;
assign twf_12_out[476] = -91;
assign twf_12_out[477] = -126;
assign twf_12_out[478] = -118;
assign twf_12_out[479] = -71;
assign twf_12_out[480] = 128;
assign twf_12_out[481] = 127;
assign twf_12_out[482] = 126;
assign twf_12_out[483] = 122;
assign twf_12_out[484] = 118;
assign twf_12_out[485] = 113;
assign twf_12_out[486] = 106;
assign twf_12_out[487] = 99;
assign twf_12_out[488] = 128;
assign twf_12_out[489] = 113;
assign twf_12_out[490] = 71;
assign twf_12_out[491] = 13;
assign twf_12_out[492] = -49;
assign twf_12_out[493] = -99;
assign twf_12_out[494] = -126;
assign twf_12_out[495] = -122;
assign twf_12_out[496] = 128;
assign twf_12_out[497] = 122;
assign twf_12_out[498] = 106;
assign twf_12_out[499] = 81;
assign twf_12_out[500] = 49;
assign twf_12_out[501] = 13;
assign twf_12_out[502] = -25;
assign twf_12_out[503] = -60;
assign twf_12_out[504] = 128;
assign twf_12_out[505] = 99;
assign twf_12_out[506] = 25;
assign twf_12_out[507] = -60;
assign twf_12_out[508] = -118;
assign twf_12_out[509] = -122;
assign twf_12_out[510] = -71;
assign twf_12_out[511] = 13;


endmodule
`timescale 1ns/1ps

module twf_12_imag #(
    parameter INDEX_WIDTH = 64,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output signed [BIT_WIDTH-1:0] twf_out
);

wire signed [BIT_WIDTH-1:0] twf_12_out [0:INDEX_WIDTH-1];

assign twf_out = twf_12_out[index];

assign twf_12_out[0] = 0;
assign twf_12_out[1] = 0;
assign twf_12_out[2] = 0;
assign twf_12_out[3] = 0;
assign twf_12_out[4] = 0;
assign twf_12_out[5] = 0;
assign twf_12_out[6] = 0;
assign twf_12_out[7] = 0;
assign twf_12_out[8] = 0;
assign twf_12_out[9] = -49;
assign twf_12_out[10] = -91;
assign twf_12_out[11] = -118;
assign twf_12_out[12] = -128;
assign twf_12_out[13] = -118;
assign twf_12_out[14] = -91;
assign twf_12_out[15] = -49;
assign twf_12_out[16] = 0;
assign twf_12_out[17] = -25;
assign twf_12_out[18] = -49;
assign twf_12_out[19] = -71;
assign twf_12_out[20] = -91;
assign twf_12_out[21] = -106;
assign twf_12_out[22] = -118;
assign twf_12_out[23] = -126;
assign twf_12_out[24] = 0;
assign twf_12_out[25] = -71;
assign twf_12_out[26] = -118;
assign twf_12_out[27] = -126;
assign twf_12_out[28] = -91;
assign twf_12_out[29] = -25;
assign twf_12_out[30] = 49;
assign twf_12_out[31] = 106;
assign twf_12_out[32] = 0;
assign twf_12_out[33] = -13;
assign twf_12_out[34] = -25;
assign twf_12_out[35] = -37;
assign twf_12_out[36] = -49;
assign twf_12_out[37] = -60;
assign twf_12_out[38] = -71;
assign twf_12_out[39] = -81;
assign twf_12_out[40] = 0;
assign twf_12_out[41] = -60;
assign twf_12_out[42] = -106;
assign twf_12_out[43] = -127;
assign twf_12_out[44] = -118;
assign twf_12_out[45] = -81;
assign twf_12_out[46] = -25;
assign twf_12_out[47] = 37;
assign twf_12_out[48] = 0;
assign twf_12_out[49] = -37;
assign twf_12_out[50] = -71;
assign twf_12_out[51] = -99;
assign twf_12_out[52] = -118;
assign twf_12_out[53] = -127;
assign twf_12_out[54] = -126;
assign twf_12_out[55] = -113;
assign twf_12_out[56] = 0;
assign twf_12_out[57] = -81;
assign twf_12_out[58] = -126;
assign twf_12_out[59] = -113;
assign twf_12_out[60] = -49;
assign twf_12_out[61] = 37;
assign twf_12_out[62] = 106;
assign twf_12_out[63] = 127;
assign twf_12_out[64] = 0;
assign twf_12_out[65] = 0;
assign twf_12_out[66] = 0;
assign twf_12_out[67] = 0;
assign twf_12_out[68] = 0;
assign twf_12_out[69] = 0;
assign twf_12_out[70] = 0;
assign twf_12_out[71] = 0;
assign twf_12_out[72] = 0;
assign twf_12_out[73] = -49;
assign twf_12_out[74] = -91;
assign twf_12_out[75] = -118;
assign twf_12_out[76] = -128;
assign twf_12_out[77] = -118;
assign twf_12_out[78] = -91;
assign twf_12_out[79] = -49;
assign twf_12_out[80] = 0;
assign twf_12_out[81] = -25;
assign twf_12_out[82] = -49;
assign twf_12_out[83] = -71;
assign twf_12_out[84] = -91;
assign twf_12_out[85] = -106;
assign twf_12_out[86] = -118;
assign twf_12_out[87] = -126;
assign twf_12_out[88] = 0;
assign twf_12_out[89] = -71;
assign twf_12_out[90] = -118;
assign twf_12_out[91] = -126;
assign twf_12_out[92] = -91;
assign twf_12_out[93] = -25;
assign twf_12_out[94] = 49;
assign twf_12_out[95] = 106;
assign twf_12_out[96] = 0;
assign twf_12_out[97] = -13;
assign twf_12_out[98] = -25;
assign twf_12_out[99] = -37;
assign twf_12_out[100] = -49;
assign twf_12_out[101] = -60;
assign twf_12_out[102] = -71;
assign twf_12_out[103] = -81;
assign twf_12_out[104] = 0;
assign twf_12_out[105] = -60;
assign twf_12_out[106] = -106;
assign twf_12_out[107] = -127;
assign twf_12_out[108] = -118;
assign twf_12_out[109] = -81;
assign twf_12_out[110] = -25;
assign twf_12_out[111] = 37;
assign twf_12_out[112] = 0;
assign twf_12_out[113] = -37;
assign twf_12_out[114] = -71;
assign twf_12_out[115] = -99;
assign twf_12_out[116] = -118;
assign twf_12_out[117] = -127;
assign twf_12_out[118] = -126;
assign twf_12_out[119] = -113;
assign twf_12_out[120] = 0;
assign twf_12_out[121] = -81;
assign twf_12_out[122] = -126;
assign twf_12_out[123] = -113;
assign twf_12_out[124] = -49;
assign twf_12_out[125] = 37;
assign twf_12_out[126] = 106;
assign twf_12_out[127] = 127;
assign twf_12_out[128] = 0;
assign twf_12_out[129] = 0;
assign twf_12_out[130] = 0;
assign twf_12_out[131] = 0;
assign twf_12_out[132] = 0;
assign twf_12_out[133] = 0;
assign twf_12_out[134] = 0;
assign twf_12_out[135] = 0;
assign twf_12_out[136] = 0;
assign twf_12_out[137] = -49;
assign twf_12_out[138] = -91;
assign twf_12_out[139] = -118;
assign twf_12_out[140] = -128;
assign twf_12_out[141] = -118;
assign twf_12_out[142] = -91;
assign twf_12_out[143] = -49;
assign twf_12_out[144] = 0;
assign twf_12_out[145] = -25;
assign twf_12_out[146] = -49;
assign twf_12_out[147] = -71;
assign twf_12_out[148] = -91;
assign twf_12_out[149] = -106;
assign twf_12_out[150] = -118;
assign twf_12_out[151] = -126;
assign twf_12_out[152] = 0;
assign twf_12_out[153] = -71;
assign twf_12_out[154] = -118;
assign twf_12_out[155] = -126;
assign twf_12_out[156] = -91;
assign twf_12_out[157] = -25;
assign twf_12_out[158] = 49;
assign twf_12_out[159] = 106;
assign twf_12_out[160] = 0;
assign twf_12_out[161] = -13;
assign twf_12_out[162] = -25;
assign twf_12_out[163] = -37;
assign twf_12_out[164] = -49;
assign twf_12_out[165] = -60;
assign twf_12_out[166] = -71;
assign twf_12_out[167] = -81;
assign twf_12_out[168] = 0;
assign twf_12_out[169] = -60;
assign twf_12_out[170] = -106;
assign twf_12_out[171] = -127;
assign twf_12_out[172] = -118;
assign twf_12_out[173] = -81;
assign twf_12_out[174] = -25;
assign twf_12_out[175] = 37;
assign twf_12_out[176] = 0;
assign twf_12_out[177] = -37;
assign twf_12_out[178] = -71;
assign twf_12_out[179] = -99;
assign twf_12_out[180] = -118;
assign twf_12_out[181] = -127;
assign twf_12_out[182] = -126;
assign twf_12_out[183] = -113;
assign twf_12_out[184] = 0;
assign twf_12_out[185] = -81;
assign twf_12_out[186] = -126;
assign twf_12_out[187] = -113;
assign twf_12_out[188] = -49;
assign twf_12_out[189] = 37;
assign twf_12_out[190] = 106;
assign twf_12_out[191] = 127;
assign twf_12_out[192] = 0;
assign twf_12_out[193] = 0;
assign twf_12_out[194] = 0;
assign twf_12_out[195] = 0;
assign twf_12_out[196] = 0;
assign twf_12_out[197] = 0;
assign twf_12_out[198] = 0;
assign twf_12_out[199] = 0;
assign twf_12_out[200] = 0;
assign twf_12_out[201] = -49;
assign twf_12_out[202] = -91;
assign twf_12_out[203] = -118;
assign twf_12_out[204] = -128;
assign twf_12_out[205] = -118;
assign twf_12_out[206] = -91;
assign twf_12_out[207] = -49;
assign twf_12_out[208] = 0;
assign twf_12_out[209] = -25;
assign twf_12_out[210] = -49;
assign twf_12_out[211] = -71;
assign twf_12_out[212] = -91;
assign twf_12_out[213] = -106;
assign twf_12_out[214] = -118;
assign twf_12_out[215] = -126;
assign twf_12_out[216] = 0;
assign twf_12_out[217] = -71;
assign twf_12_out[218] = -118;
assign twf_12_out[219] = -126;
assign twf_12_out[220] = -91;
assign twf_12_out[221] = -25;
assign twf_12_out[222] = 49;
assign twf_12_out[223] = 106;
assign twf_12_out[224] = 0;
assign twf_12_out[225] = -13;
assign twf_12_out[226] = -25;
assign twf_12_out[227] = -37;
assign twf_12_out[228] = -49;
assign twf_12_out[229] = -60;
assign twf_12_out[230] = -71;
assign twf_12_out[231] = -81;
assign twf_12_out[232] = 0;
assign twf_12_out[233] = -60;
assign twf_12_out[234] = -106;
assign twf_12_out[235] = -127;
assign twf_12_out[236] = -118;
assign twf_12_out[237] = -81;
assign twf_12_out[238] = -25;
assign twf_12_out[239] = 37;
assign twf_12_out[240] = 0;
assign twf_12_out[241] = -37;
assign twf_12_out[242] = -71;
assign twf_12_out[243] = -99;
assign twf_12_out[244] = -118;
assign twf_12_out[245] = -127;
assign twf_12_out[246] = -126;
assign twf_12_out[247] = -113;
assign twf_12_out[248] = 0;
assign twf_12_out[249] = -81;
assign twf_12_out[250] = -126;
assign twf_12_out[251] = -113;
assign twf_12_out[252] = -49;
assign twf_12_out[253] = 37;
assign twf_12_out[254] = 106;
assign twf_12_out[255] = 127;
assign twf_12_out[256] = 0;
assign twf_12_out[257] = 0;
assign twf_12_out[258] = 0;
assign twf_12_out[259] = 0;
assign twf_12_out[260] = 0;
assign twf_12_out[261] = 0;
assign twf_12_out[262] = 0;
assign twf_12_out[263] = 0;
assign twf_12_out[264] = 0;
assign twf_12_out[265] = -49;
assign twf_12_out[266] = -91;
assign twf_12_out[267] = -118;
assign twf_12_out[268] = -128;
assign twf_12_out[269] = -118;
assign twf_12_out[270] = -91;
assign twf_12_out[271] = -49;
assign twf_12_out[272] = 0;
assign twf_12_out[273] = -25;
assign twf_12_out[274] = -49;
assign twf_12_out[275] = -71;
assign twf_12_out[276] = -91;
assign twf_12_out[277] = -106;
assign twf_12_out[278] = -118;
assign twf_12_out[279] = -126;
assign twf_12_out[280] = 0;
assign twf_12_out[281] = -71;
assign twf_12_out[282] = -118;
assign twf_12_out[283] = -126;
assign twf_12_out[284] = -91;
assign twf_12_out[285] = -25;
assign twf_12_out[286] = 49;
assign twf_12_out[287] = 106;
assign twf_12_out[288] = 0;
assign twf_12_out[289] = -13;
assign twf_12_out[290] = -25;
assign twf_12_out[291] = -37;
assign twf_12_out[292] = -49;
assign twf_12_out[293] = -60;
assign twf_12_out[294] = -71;
assign twf_12_out[295] = -81;
assign twf_12_out[296] = 0;
assign twf_12_out[297] = -60;
assign twf_12_out[298] = -106;
assign twf_12_out[299] = -127;
assign twf_12_out[300] = -118;
assign twf_12_out[301] = -81;
assign twf_12_out[302] = -25;
assign twf_12_out[303] = 37;
assign twf_12_out[304] = 0;
assign twf_12_out[305] = -37;
assign twf_12_out[306] = -71;
assign twf_12_out[307] = -99;
assign twf_12_out[308] = -118;
assign twf_12_out[309] = -127;
assign twf_12_out[310] = -126;
assign twf_12_out[311] = -113;
assign twf_12_out[312] = 0;
assign twf_12_out[313] = -81;
assign twf_12_out[314] = -126;
assign twf_12_out[315] = -113;
assign twf_12_out[316] = -49;
assign twf_12_out[317] = 37;
assign twf_12_out[318] = 106;
assign twf_12_out[319] = 127;
assign twf_12_out[320] = 0;
assign twf_12_out[321] = 0;
assign twf_12_out[322] = 0;
assign twf_12_out[323] = 0;
assign twf_12_out[324] = 0;
assign twf_12_out[325] = 0;
assign twf_12_out[326] = 0;
assign twf_12_out[327] = 0;
assign twf_12_out[328] = 0;
assign twf_12_out[329] = -49;
assign twf_12_out[330] = -91;
assign twf_12_out[331] = -118;
assign twf_12_out[332] = -128;
assign twf_12_out[333] = -118;
assign twf_12_out[334] = -91;
assign twf_12_out[335] = -49;
assign twf_12_out[336] = 0;
assign twf_12_out[337] = -25;
assign twf_12_out[338] = -49;
assign twf_12_out[339] = -71;
assign twf_12_out[340] = -91;
assign twf_12_out[341] = -106;
assign twf_12_out[342] = -118;
assign twf_12_out[343] = -126;
assign twf_12_out[344] = 0;
assign twf_12_out[345] = -71;
assign twf_12_out[346] = -118;
assign twf_12_out[347] = -126;
assign twf_12_out[348] = -91;
assign twf_12_out[349] = -25;
assign twf_12_out[350] = 49;
assign twf_12_out[351] = 106;
assign twf_12_out[352] = 0;
assign twf_12_out[353] = -13;
assign twf_12_out[354] = -25;
assign twf_12_out[355] = -37;
assign twf_12_out[356] = -49;
assign twf_12_out[357] = -60;
assign twf_12_out[358] = -71;
assign twf_12_out[359] = -81;
assign twf_12_out[360] = 0;
assign twf_12_out[361] = -60;
assign twf_12_out[362] = -106;
assign twf_12_out[363] = -127;
assign twf_12_out[364] = -118;
assign twf_12_out[365] = -81;
assign twf_12_out[366] = -25;
assign twf_12_out[367] = 37;
assign twf_12_out[368] = 0;
assign twf_12_out[369] = -37;
assign twf_12_out[370] = -71;
assign twf_12_out[371] = -99;
assign twf_12_out[372] = -118;
assign twf_12_out[373] = -127;
assign twf_12_out[374] = -126;
assign twf_12_out[375] = -113;
assign twf_12_out[376] = 0;
assign twf_12_out[377] = -81;
assign twf_12_out[378] = -126;
assign twf_12_out[379] = -113;
assign twf_12_out[380] = -49;
assign twf_12_out[381] = 37;
assign twf_12_out[382] = 106;
assign twf_12_out[383] = 127;
assign twf_12_out[384] = 0;
assign twf_12_out[385] = 0;
assign twf_12_out[386] = 0;
assign twf_12_out[387] = 0;
assign twf_12_out[388] = 0;
assign twf_12_out[389] = 0;
assign twf_12_out[390] = 0;
assign twf_12_out[391] = 0;
assign twf_12_out[392] = 0;
assign twf_12_out[393] = -49;
assign twf_12_out[394] = -91;
assign twf_12_out[395] = -118;
assign twf_12_out[396] = -128;
assign twf_12_out[397] = -118;
assign twf_12_out[398] = -91;
assign twf_12_out[399] = -49;
assign twf_12_out[400] = 0;
assign twf_12_out[401] = -25;
assign twf_12_out[402] = -49;
assign twf_12_out[403] = -71;
assign twf_12_out[404] = -91;
assign twf_12_out[405] = -106;
assign twf_12_out[406] = -118;
assign twf_12_out[407] = -126;
assign twf_12_out[408] = 0;
assign twf_12_out[409] = -71;
assign twf_12_out[410] = -118;
assign twf_12_out[411] = -126;
assign twf_12_out[412] = -91;
assign twf_12_out[413] = -25;
assign twf_12_out[414] = 49;
assign twf_12_out[415] = 106;
assign twf_12_out[416] = 0;
assign twf_12_out[417] = -13;
assign twf_12_out[418] = -25;
assign twf_12_out[419] = -37;
assign twf_12_out[420] = -49;
assign twf_12_out[421] = -60;
assign twf_12_out[422] = -71;
assign twf_12_out[423] = -81;
assign twf_12_out[424] = 0;
assign twf_12_out[425] = -60;
assign twf_12_out[426] = -106;
assign twf_12_out[427] = -127;
assign twf_12_out[428] = -118;
assign twf_12_out[429] = -81;
assign twf_12_out[430] = -25;
assign twf_12_out[431] = 37;
assign twf_12_out[432] = 0;
assign twf_12_out[433] = -37;
assign twf_12_out[434] = -71;
assign twf_12_out[435] = -99;
assign twf_12_out[436] = -118;
assign twf_12_out[437] = -127;
assign twf_12_out[438] = -126;
assign twf_12_out[439] = -113;
assign twf_12_out[440] = 0;
assign twf_12_out[441] = -81;
assign twf_12_out[442] = -126;
assign twf_12_out[443] = -113;
assign twf_12_out[444] = -49;
assign twf_12_out[445] = 37;
assign twf_12_out[446] = 106;
assign twf_12_out[447] = 127;
assign twf_12_out[448] = 0;
assign twf_12_out[449] = 0;
assign twf_12_out[450] = 0;
assign twf_12_out[451] = 0;
assign twf_12_out[452] = 0;
assign twf_12_out[453] = 0;
assign twf_12_out[454] = 0;
assign twf_12_out[455] = 0;
assign twf_12_out[456] = 0;
assign twf_12_out[457] = -49;
assign twf_12_out[458] = -91;
assign twf_12_out[459] = -118;
assign twf_12_out[460] = -128;
assign twf_12_out[461] = -118;
assign twf_12_out[462] = -91;
assign twf_12_out[463] = -49;
assign twf_12_out[464] = 0;
assign twf_12_out[465] = -25;
assign twf_12_out[466] = -49;
assign twf_12_out[467] = -71;
assign twf_12_out[468] = -91;
assign twf_12_out[469] = -106;
assign twf_12_out[470] = -118;
assign twf_12_out[471] = -126;
assign twf_12_out[472] = 0;
assign twf_12_out[473] = -71;
assign twf_12_out[474] = -118;
assign twf_12_out[475] = -126;
assign twf_12_out[476] = -91;
assign twf_12_out[477] = -25;
assign twf_12_out[478] = 49;
assign twf_12_out[479] = 106;
assign twf_12_out[480] = 0;
assign twf_12_out[481] = -13;
assign twf_12_out[482] = -25;
assign twf_12_out[483] = -37;
assign twf_12_out[484] = -49;
assign twf_12_out[485] = -60;
assign twf_12_out[486] = -71;
assign twf_12_out[487] = -81;
assign twf_12_out[488] = 0;
assign twf_12_out[489] = -60;
assign twf_12_out[490] = -106;
assign twf_12_out[491] = -127;
assign twf_12_out[492] = -118;
assign twf_12_out[493] = -81;
assign twf_12_out[494] = -25;
assign twf_12_out[495] = 37;
assign twf_12_out[496] = 0;
assign twf_12_out[497] = -37;
assign twf_12_out[498] = -71;
assign twf_12_out[499] = -99;
assign twf_12_out[500] = -118;
assign twf_12_out[501] = -127;
assign twf_12_out[502] = -126;
assign twf_12_out[503] = -113;
assign twf_12_out[504] = 0;
assign twf_12_out[505] = -81;
assign twf_12_out[506] = -126;
assign twf_12_out[507] = -113;
assign twf_12_out[508] = -49;
assign twf_12_out[509] = 37;
assign twf_12_out[510] = 106;
assign twf_12_out[511] = 127;

endmodule
module shifter #(
    parameters N = 12;
) (
    
);
    
endmodule
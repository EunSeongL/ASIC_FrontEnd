`timescale 1ns/1ps

module twf_12_imag #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output logic signed [BIT_WIDTH-1:0] twf_out
);

always @(*) begin
    case(index)
        0: twf_out = 0;
        1: twf_out = 0;
        2: twf_out = 0;
        3: twf_out = 0;
        4: twf_out = 0;
        5: twf_out = 0;
        6: twf_out = 0;
        7: twf_out = 0;
        8: twf_out = 0;
        9: twf_out = -49;
        10: twf_out = -91;
        11: twf_out = -118;
        12: twf_out = -128;
        13: twf_out = -118;
        14: twf_out = -91;
        15: twf_out = -49;
        16: twf_out = 0;
        17: twf_out = -25;
        18: twf_out = -49;
        19: twf_out = -71;
        20: twf_out = -91;
        21: twf_out = -106;
        22: twf_out = -118;
        23: twf_out = -126;
        24: twf_out = 0;
        25: twf_out = -71;
        26: twf_out = -118;
        27: twf_out = -126;
        28: twf_out = -91;
        29: twf_out = -25;
        30: twf_out = 49;
        31: twf_out = 106;
        32: twf_out = 0;
        33: twf_out = -13;
        34: twf_out = -25;
        35: twf_out = -37;
        36: twf_out = -49;
        37: twf_out = -60;
        38: twf_out = -71;
        39: twf_out = -81;
        40: twf_out = 0;
        41: twf_out = -60;
        42: twf_out = -106;
        43: twf_out = -127;
        44: twf_out = -118;
        45: twf_out = -81;
        46: twf_out = -25;
        47: twf_out = 37;
        48: twf_out = 0;
        49: twf_out = -37;
        50: twf_out = -71;
        51: twf_out = -99;
        52: twf_out = -118;
        53: twf_out = -127;
        54: twf_out = -126;
        55: twf_out = -113;
        56: twf_out = 0;
        57: twf_out = -81;
        58: twf_out = -126;
        59: twf_out = -113;
        60: twf_out = -49;
        61: twf_out = 37;
        62: twf_out = 106;
        63: twf_out = 127;
        64: twf_out = 0;
        65: twf_out = 0;
        66: twf_out = 0;
        67: twf_out = 0;
        68: twf_out = 0;
        69: twf_out = 0;
        70: twf_out = 0;
        71: twf_out = 0;
        72: twf_out = 0;
        73: twf_out = -49;
        74: twf_out = -91;
        75: twf_out = -118;
        76: twf_out = -128;
        77: twf_out = -118;
        78: twf_out = -91;
        79: twf_out = -49;
        80: twf_out = 0;
        81: twf_out = -25;
        82: twf_out = -49;
        83: twf_out = -71;
        84: twf_out = -91;
        85: twf_out = -106;
        86: twf_out = -118;
        87: twf_out = -126;
        88: twf_out = 0;
        89: twf_out = -71;
        90: twf_out = -118;
        91: twf_out = -126;
        92: twf_out = -91;
        93: twf_out = -25;
        94: twf_out = 49;
        95: twf_out = 106;
        96: twf_out = 0;
        97: twf_out = -13;
        98: twf_out = -25;
        99: twf_out = -37;
        100: twf_out = -49;
        101: twf_out = -60;
        102: twf_out = -71;
        103: twf_out = -81;
        104: twf_out = 0;
        105: twf_out = -60;
        106: twf_out = -106;
        107: twf_out = -127;
        108: twf_out = -118;
        109: twf_out = -81;
        110: twf_out = -25;
        111: twf_out = 37;
        112: twf_out = 0;
        113: twf_out = -37;
        114: twf_out = -71;
        115: twf_out = -99;
        116: twf_out = -118;
        117: twf_out = -127;
        118: twf_out = -126;
        119: twf_out = -113;
        120: twf_out = 0;
        121: twf_out = -81;
        122: twf_out = -126;
        123: twf_out = -113;
        124: twf_out = -49;
        125: twf_out = 37;
        126: twf_out = 106;
        127: twf_out = 127;
        128: twf_out = 0;
        129: twf_out = 0;
        130: twf_out = 0;
        131: twf_out = 0;
        132: twf_out = 0;
        133: twf_out = 0;
        134: twf_out = 0;
        135: twf_out = 0;
        136: twf_out = 0;
        137: twf_out = -49;
        138: twf_out = -91;
        139: twf_out = -118;
        140: twf_out = -128;
        141: twf_out = -118;
        142: twf_out = -91;
        143: twf_out = -49;
        144: twf_out = 0;
        145: twf_out = -25;
        146: twf_out = -49;
        147: twf_out = -71;
        148: twf_out = -91;
        149: twf_out = -106;
        150: twf_out = -118;
        151: twf_out = -126;
        152: twf_out = 0;
        153: twf_out = -71;
        154: twf_out = -118;
        155: twf_out = -126;
        156: twf_out = -91;
        157: twf_out = -25;
        158: twf_out = 49;
        159: twf_out = 106;
        160: twf_out = 0;
        161: twf_out = -13;
        162: twf_out = -25;
        163: twf_out = -37;
        164: twf_out = -49;
        165: twf_out = -60;
        166: twf_out = -71;
        167: twf_out = -81;
        168: twf_out = 0;
        169: twf_out = -60;
        170: twf_out = -106;
        171: twf_out = -127;
        172: twf_out = -118;
        173: twf_out = -81;
        174: twf_out = -25;
        175: twf_out = 37;
        176: twf_out = 0;
        177: twf_out = -37;
        178: twf_out = -71;
        179: twf_out = -99;
        180: twf_out = -118;
        181: twf_out = -127;
        182: twf_out = -126;
        183: twf_out = -113;
        184: twf_out = 0;
        185: twf_out = -81;
        186: twf_out = -126;
        187: twf_out = -113;
        188: twf_out = -49;
        189: twf_out = 37;
        190: twf_out = 106;
        191: twf_out = 127;
        192: twf_out = 0;
        193: twf_out = 0;
        194: twf_out = 0;
        195: twf_out = 0;
        196: twf_out = 0;
        197: twf_out = 0;
        198: twf_out = 0;
        199: twf_out = 0;
        200: twf_out = 0;
        201: twf_out = -49;
        202: twf_out = -91;
        203: twf_out = -118;
        204: twf_out = -128;
        205: twf_out = -118;
        206: twf_out = -91;
        207: twf_out = -49;
        208: twf_out = 0;
        209: twf_out = -25;
        210: twf_out = -49;
        211: twf_out = -71;
        212: twf_out = -91;
        213: twf_out = -106;
        214: twf_out = -118;
        215: twf_out = -126;
        216: twf_out = 0;
        217: twf_out = -71;
        218: twf_out = -118;
        219: twf_out = -126;
        220: twf_out = -91;
        221: twf_out = -25;
        222: twf_out = 49;
        223: twf_out = 106;
        224: twf_out = 0;
        225: twf_out = -13;
        226: twf_out = -25;
        227: twf_out = -37;
        228: twf_out = -49;
        229: twf_out = -60;
        230: twf_out = -71;
        231: twf_out = -81;
        232: twf_out = 0;
        233: twf_out = -60;
        234: twf_out = -106;
        235: twf_out = -127;
        236: twf_out = -118;
        237: twf_out = -81;
        238: twf_out = -25;
        239: twf_out = 37;
        240: twf_out = 0;
        241: twf_out = -37;
        242: twf_out = -71;
        243: twf_out = -99;
        244: twf_out = -118;
        245: twf_out = -127;
        246: twf_out = -126;
        247: twf_out = -113;
        248: twf_out = 0;
        249: twf_out = -81;
        250: twf_out = -126;
        251: twf_out = -113;
        252: twf_out = -49;
        253: twf_out = 37;
        254: twf_out = 106;
        255: twf_out = 127;
        256: twf_out = 0;
        257: twf_out = 0;
        258: twf_out = 0;
        259: twf_out = 0;
        260: twf_out = 0;
        261: twf_out = 0;
        262: twf_out = 0;
        263: twf_out = 0;
        264: twf_out = 0;
        265: twf_out = -49;
        266: twf_out = -91;
        267: twf_out = -118;
        268: twf_out = -128;
        269: twf_out = -118;
        270: twf_out = -91;
        271: twf_out = -49;
        272: twf_out = 0;
        273: twf_out = -25;
        274: twf_out = -49;
        275: twf_out = -71;
        276: twf_out = -91;
        277: twf_out = -106;
        278: twf_out = -118;
        279: twf_out = -126;
        280: twf_out = 0;
        281: twf_out = -71;
        282: twf_out = -118;
        283: twf_out = -126;
        284: twf_out = -91;
        285: twf_out = -25;
        286: twf_out = 49;
        287: twf_out = 106;
        288: twf_out = 0;
        289: twf_out = -13;
        290: twf_out = -25;
        291: twf_out = -37;
        292: twf_out = -49;
        293: twf_out = -60;
        294: twf_out = -71;
        295: twf_out = -81;
        296: twf_out = 0;
        297: twf_out = -60;
        298: twf_out = -106;
        299: twf_out = -127;
        300: twf_out = -118;
        301: twf_out = -81;
        302: twf_out = -25;
        303: twf_out = 37;
        304: twf_out = 0;
        305: twf_out = -37;
        306: twf_out = -71;
        307: twf_out = -99;
        308: twf_out = -118;
        309: twf_out = -127;
        310: twf_out = -126;
        311: twf_out = -113;
        312: twf_out = 0;
        313: twf_out = -81;
        314: twf_out = -126;
        315: twf_out = -113;
        316: twf_out = -49;
        317: twf_out = 37;
        318: twf_out = 106;
        319: twf_out = 127;
        320: twf_out = 0;
        321: twf_out = 0;
        322: twf_out = 0;
        323: twf_out = 0;
        324: twf_out = 0;
        325: twf_out = 0;
        326: twf_out = 0;
        327: twf_out = 0;
        328: twf_out = 0;
        329: twf_out = -49;
        330: twf_out = -91;
        331: twf_out = -118;
        332: twf_out = -128;
        333: twf_out = -118;
        334: twf_out = -91;
        335: twf_out = -49;
        336: twf_out = 0;
        337: twf_out = -25;
        338: twf_out = -49;
        339: twf_out = -71;
        340: twf_out = -91;
        341: twf_out = -106;
        342: twf_out = -118;
        343: twf_out = -126;
        344: twf_out = 0;
        345: twf_out = -71;
        346: twf_out = -118;
        347: twf_out = -126;
        348: twf_out = -91;
        349: twf_out = -25;
        350: twf_out = 49;
        351: twf_out = 106;
        352: twf_out = 0;
        353: twf_out = -13;
        354: twf_out = -25;
        355: twf_out = -37;
        356: twf_out = -49;
        357: twf_out = -60;
        358: twf_out = -71;
        359: twf_out = -81;
        360: twf_out = 0;
        361: twf_out = -60;
        362: twf_out = -106;
        363: twf_out = -127;
        364: twf_out = -118;
        365: twf_out = -81;
        366: twf_out = -25;
        367: twf_out = 37;
        368: twf_out = 0;
        369: twf_out = -37;
        370: twf_out = -71;
        371: twf_out = -99;
        372: twf_out = -118;
        373: twf_out = -127;
        374: twf_out = -126;
        375: twf_out = -113;
        376: twf_out = 0;
        377: twf_out = -81;
        378: twf_out = -126;
        379: twf_out = -113;
        380: twf_out = -49;
        381: twf_out = 37;
        382: twf_out = 106;
        383: twf_out = 127;
        384: twf_out = 0;
        385: twf_out = 0;
        386: twf_out = 0;
        387: twf_out = 0;
        388: twf_out = 0;
        389: twf_out = 0;
        390: twf_out = 0;
        391: twf_out = 0;
        392: twf_out = 0;
        393: twf_out = -49;
        394: twf_out = -91;
        395: twf_out = -118;
        396: twf_out = -128;
        397: twf_out = -118;
        398: twf_out = -91;
        399: twf_out = -49;
        400: twf_out = 0;
        401: twf_out = -25;
        402: twf_out = -49;
        403: twf_out = -71;
        404: twf_out = -91;
        405: twf_out = -106;
        406: twf_out = -118;
        407: twf_out = -126;
        408: twf_out = 0;
        409: twf_out = -71;
        410: twf_out = -118;
        411: twf_out = -126;
        412: twf_out = -91;
        413: twf_out = -25;
        414: twf_out = 49;
        415: twf_out = 106;
        416: twf_out = 0;
        417: twf_out = -13;
        418: twf_out = -25;
        419: twf_out = -37;
        420: twf_out = -49;
        421: twf_out = -60;
        422: twf_out = -71;
        423: twf_out = -81;
        424: twf_out = 0;
        425: twf_out = -60;
        426: twf_out = -106;
        427: twf_out = -127;
        428: twf_out = -118;
        429: twf_out = -81;
        430: twf_out = -25;
        431: twf_out = 37;
        432: twf_out = 0;
        433: twf_out = -37;
        434: twf_out = -71;
        435: twf_out = -99;
        436: twf_out = -118;
        437: twf_out = -127;
        438: twf_out = -126;
        439: twf_out = -113;
        440: twf_out = 0;
        441: twf_out = -81;
        442: twf_out = -126;
        443: twf_out = -113;
        444: twf_out = -49;
        445: twf_out = 37;
        446: twf_out = 106;
        447: twf_out = 127;
        448: twf_out = 0;
        449: twf_out = 0;
        450: twf_out = 0;
        451: twf_out = 0;
        452: twf_out = 0;
        453: twf_out = 0;
        454: twf_out = 0;
        455: twf_out = 0;
        456: twf_out = 0;
        457: twf_out = -49;
        458: twf_out = -91;
        459: twf_out = -118;
        460: twf_out = -128;
        461: twf_out = -118;
        462: twf_out = -91;
        463: twf_out = -49;
        464: twf_out = 0;
        465: twf_out = -25;
        466: twf_out = -49;
        467: twf_out = -71;
        468: twf_out = -91;
        469: twf_out = -106;
        470: twf_out = -118;
        471: twf_out = -126;
        472: twf_out = 0;
        473: twf_out = -71;
        474: twf_out = -118;
        475: twf_out = -126;
        476: twf_out = -91;
        477: twf_out = -25;
        478: twf_out = 49;
        479: twf_out = 106;
        480: twf_out = 0;
        481: twf_out = -13;
        482: twf_out = -25;
        483: twf_out = -37;
        484: twf_out = -49;
        485: twf_out = -60;
        486: twf_out = -71;
        487: twf_out = -81;
        488: twf_out = 0;
        489: twf_out = -60;
        490: twf_out = -106;
        491: twf_out = -127;
        492: twf_out = -118;
        493: twf_out = -81;
        494: twf_out = -25;
        495: twf_out = 37;
        496: twf_out = 0;
        497: twf_out = -37;
        498: twf_out = -71;
        499: twf_out = -99;
        500: twf_out = -118;
        501: twf_out = -127;
        502: twf_out = -126;
        503: twf_out = -113;
        504: twf_out = 0;
        505: twf_out = -81;
        506: twf_out = -126;
        507: twf_out = -113;
        508: twf_out = -49;
        509: twf_out = 37;
        510: twf_out = 106;
        511: twf_out = 127;
        default: twf_out = 0;
    endcase
end

endmodule

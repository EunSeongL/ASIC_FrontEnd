`timescale 1ns/1ps

module twf_12_real #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output logic signed [BIT_WIDTH-1:0] twf_out
);

always @(*) begin
    case(index)
        0: twf_out = 128;
        1: twf_out = 128;
        2: twf_out = 128;
        3: twf_out = 128;
        4: twf_out = 128;
        5: twf_out = 128;
        6: twf_out = 128;
        7: twf_out = 128;
        8: twf_out = 128;
        9: twf_out = 118;
        10: twf_out = 91;
        11: twf_out = 49;
        12: twf_out = 0;
        13: twf_out = -49;
        14: twf_out = -91;
        15: twf_out = -118;
        16: twf_out = 128;
        17: twf_out = 126;
        18: twf_out = 118;
        19: twf_out = 106;
        20: twf_out = 91;
        21: twf_out = 71;
        22: twf_out = 49;
        23: twf_out = 25;
        24: twf_out = 128;
        25: twf_out = 106;
        26: twf_out = 49;
        27: twf_out = -25;
        28: twf_out = -91;
        29: twf_out = -126;
        30: twf_out = -118;
        31: twf_out = -71;
        32: twf_out = 128;
        33: twf_out = 127;
        34: twf_out = 126;
        35: twf_out = 122;
        36: twf_out = 118;
        37: twf_out = 113;
        38: twf_out = 106;
        39: twf_out = 99;
        40: twf_out = 128;
        41: twf_out = 113;
        42: twf_out = 71;
        43: twf_out = 13;
        44: twf_out = -49;
        45: twf_out = -99;
        46: twf_out = -126;
        47: twf_out = -122;
        48: twf_out = 128;
        49: twf_out = 122;
        50: twf_out = 106;
        51: twf_out = 81;
        52: twf_out = 49;
        53: twf_out = 13;
        54: twf_out = -25;
        55: twf_out = -60;
        56: twf_out = 128;
        57: twf_out = 99;
        58: twf_out = 25;
        59: twf_out = -60;
        60: twf_out = -118;
        61: twf_out = -122;
        62: twf_out = -71;
        63: twf_out = 13;
        64: twf_out = 128;
        65: twf_out = 128;
        66: twf_out = 128;
        67: twf_out = 128;
        68: twf_out = 128;
        69: twf_out = 128;
        70: twf_out = 128;
        71: twf_out = 128;
        72: twf_out = 128;
        73: twf_out = 118;
        74: twf_out = 91;
        75: twf_out = 49;
        76: twf_out = 0;
        77: twf_out = -49;
        78: twf_out = -91;
        79: twf_out = -118;
        80: twf_out = 128;
        81: twf_out = 126;
        82: twf_out = 118;
        83: twf_out = 106;
        84: twf_out = 91;
        85: twf_out = 71;
        86: twf_out = 49;
        87: twf_out = 25;
        88: twf_out = 128;
        89: twf_out = 106;
        90: twf_out = 49;
        91: twf_out = -25;
        92: twf_out = -91;
        93: twf_out = -126;
        94: twf_out = -118;
        95: twf_out = -71;
        96: twf_out = 128;
        97: twf_out = 127;
        98: twf_out = 126;
        99: twf_out = 122;
        100: twf_out = 118;
        101: twf_out = 113;
        102: twf_out = 106;
        103: twf_out = 99;
        104: twf_out = 128;
        105: twf_out = 113;
        106: twf_out = 71;
        107: twf_out = 13;
        108: twf_out = -49;
        109: twf_out = -99;
        110: twf_out = -126;
        111: twf_out = -122;
        112: twf_out = 128;
        113: twf_out = 122;
        114: twf_out = 106;
        115: twf_out = 81;
        116: twf_out = 49;
        117: twf_out = 13;
        118: twf_out = -25;
        119: twf_out = -60;
        120: twf_out = 128;
        121: twf_out = 99;
        122: twf_out = 25;
        123: twf_out = -60;
        124: twf_out = -118;
        125: twf_out = -122;
        126: twf_out = -71;
        127: twf_out = 13;
        128: twf_out = 128;
        129: twf_out = 128;
        130: twf_out = 128;
        131: twf_out = 128;
        132: twf_out = 128;
        133: twf_out = 128;
        134: twf_out = 128;
        135: twf_out = 128;
        136: twf_out = 128;
        137: twf_out = 118;
        138: twf_out = 91;
        139: twf_out = 49;
        140: twf_out = 0;
        141: twf_out = -49;
        142: twf_out = -91;
        143: twf_out = -118;
        144: twf_out = 128;
        145: twf_out = 126;
        146: twf_out = 118;
        147: twf_out = 106;
        148: twf_out = 91;
        149: twf_out = 71;
        150: twf_out = 49;
        151: twf_out = 25;
        152: twf_out = 128;
        153: twf_out = 106;
        154: twf_out = 49;
        155: twf_out = -25;
        156: twf_out = -91;
        157: twf_out = -126;
        158: twf_out = -118;
        159: twf_out = -71;
        160: twf_out = 128;
        161: twf_out = 127;
        162: twf_out = 126;
        163: twf_out = 122;
        164: twf_out = 118;
        165: twf_out = 113;
        166: twf_out = 106;
        167: twf_out = 99;
        168: twf_out = 128;
        169: twf_out = 113;
        170: twf_out = 71;
        171: twf_out = 13;
        172: twf_out = -49;
        173: twf_out = -99;
        174: twf_out = -126;
        175: twf_out = -122;
        176: twf_out = 128;
        177: twf_out = 122;
        178: twf_out = 106;
        179: twf_out = 81;
        180: twf_out = 49;
        181: twf_out = 13;
        182: twf_out = -25;
        183: twf_out = -60;
        184: twf_out = 128;
        185: twf_out = 99;
        186: twf_out = 25;
        187: twf_out = -60;
        188: twf_out = -118;
        189: twf_out = -122;
        190: twf_out = -71;
        191: twf_out = 13;
        192: twf_out = 128;
        193: twf_out = 128;
        194: twf_out = 128;
        195: twf_out = 128;
        196: twf_out = 128;
        197: twf_out = 128;
        198: twf_out = 128;
        199: twf_out = 128;
        200: twf_out = 128;
        201: twf_out = 118;
        202: twf_out = 91;
        203: twf_out = 49;
        204: twf_out = 0;
        205: twf_out = -49;
        206: twf_out = -91;
        207: twf_out = -118;
        208: twf_out = 128;
        209: twf_out = 126;
        210: twf_out = 118;
        211: twf_out = 106;
        212: twf_out = 91;
        213: twf_out = 71;
        214: twf_out = 49;
        215: twf_out = 25;
        216: twf_out = 128;
        217: twf_out = 106;
        218: twf_out = 49;
        219: twf_out = -25;
        220: twf_out = -91;
        221: twf_out = -126;
        222: twf_out = -118;
        223: twf_out = -71;
        224: twf_out = 128;
        225: twf_out = 127;
        226: twf_out = 126;
        227: twf_out = 122;
        228: twf_out = 118;
        229: twf_out = 113;
        230: twf_out = 106;
        231: twf_out = 99;
        232: twf_out = 128;
        233: twf_out = 113;
        234: twf_out = 71;
        235: twf_out = 13;
        236: twf_out = -49;
        237: twf_out = -99;
        238: twf_out = -126;
        239: twf_out = -122;
        240: twf_out = 128;
        241: twf_out = 122;
        242: twf_out = 106;
        243: twf_out = 81;
        244: twf_out = 49;
        245: twf_out = 13;
        246: twf_out = -25;
        247: twf_out = -60;
        248: twf_out = 128;
        249: twf_out = 99;
        250: twf_out = 25;
        251: twf_out = -60;
        252: twf_out = -118;
        253: twf_out = -122;
        254: twf_out = -71;
        255: twf_out = 13;
        256: twf_out = 128;
        257: twf_out = 128;
        258: twf_out = 128;
        259: twf_out = 128;
        260: twf_out = 128;
        261: twf_out = 128;
        262: twf_out = 128;
        263: twf_out = 128;
        264: twf_out = 128;
        265: twf_out = 118;
        266: twf_out = 91;
        267: twf_out = 49;
        268: twf_out = 0;
        269: twf_out = -49;
        270: twf_out = -91;
        271: twf_out = -118;
        272: twf_out = 128;
        273: twf_out = 126;
        274: twf_out = 118;
        275: twf_out = 106;
        276: twf_out = 91;
        277: twf_out = 71;
        278: twf_out = 49;
        279: twf_out = 25;
        280: twf_out = 128;
        281: twf_out = 106;
        282: twf_out = 49;
        283: twf_out = -25;
        284: twf_out = -91;
        285: twf_out = -126;
        286: twf_out = -118;
        287: twf_out = -71;
        288: twf_out = 128;
        289: twf_out = 127;
        290: twf_out = 126;
        291: twf_out = 122;
        292: twf_out = 118;
        293: twf_out = 113;
        294: twf_out = 106;
        295: twf_out = 99;
        296: twf_out = 128;
        297: twf_out = 113;
        298: twf_out = 71;
        299: twf_out = 13;
        300: twf_out = -49;
        301: twf_out = -99;
        302: twf_out = -126;
        303: twf_out = -122;
        304: twf_out = 128;
        305: twf_out = 122;
        306: twf_out = 106;
        307: twf_out = 81;
        308: twf_out = 49;
        309: twf_out = 13;
        310: twf_out = -25;
        311: twf_out = -60;
        312: twf_out = 128;
        313: twf_out = 99;
        314: twf_out = 25;
        315: twf_out = -60;
        316: twf_out = -118;
        317: twf_out = -122;
        318: twf_out = -71;
        319: twf_out = 13;
        320: twf_out = 128;
        321: twf_out = 128;
        322: twf_out = 128;
        323: twf_out = 128;
        324: twf_out = 128;
        325: twf_out = 128;
        326: twf_out = 128;
        327: twf_out = 128;
        328: twf_out = 128;
        329: twf_out = 118;
        330: twf_out = 91;
        331: twf_out = 49;
        332: twf_out = 0;
        333: twf_out = -49;
        334: twf_out = -91;
        335: twf_out = -118;
        336: twf_out = 128;
        337: twf_out = 126;
        338: twf_out = 118;
        339: twf_out = 106;
        340: twf_out = 91;
        341: twf_out = 71;
        342: twf_out = 49;
        343: twf_out = 25;
        344: twf_out = 128;
        345: twf_out = 106;
        346: twf_out = 49;
        347: twf_out = -25;
        348: twf_out = -91;
        349: twf_out = -126;
        350: twf_out = -118;
        351: twf_out = -71;
        352: twf_out = 128;
        353: twf_out = 127;
        354: twf_out = 126;
        355: twf_out = 122;
        356: twf_out = 118;
        357: twf_out = 113;
        358: twf_out = 106;
        359: twf_out = 99;
        360: twf_out = 128;
        361: twf_out = 113;
        362: twf_out = 71;
        363: twf_out = 13;
        364: twf_out = -49;
        365: twf_out = -99;
        366: twf_out = -126;
        367: twf_out = -122;
        368: twf_out = 128;
        369: twf_out = 122;
        370: twf_out = 106;
        371: twf_out = 81;
        372: twf_out = 49;
        373: twf_out = 13;
        374: twf_out = -25;
        375: twf_out = -60;
        376: twf_out = 128;
        377: twf_out = 99;
        378: twf_out = 25;
        379: twf_out = -60;
        380: twf_out = -118;
        381: twf_out = -122;
        382: twf_out = -71;
        383: twf_out = 13;
        384: twf_out = 128;
        385: twf_out = 128;
        386: twf_out = 128;
        387: twf_out = 128;
        388: twf_out = 128;
        389: twf_out = 128;
        390: twf_out = 128;
        391: twf_out = 128;
        392: twf_out = 128;
        393: twf_out = 118;
        394: twf_out = 91;
        395: twf_out = 49;
        396: twf_out = 0;
        397: twf_out = -49;
        398: twf_out = -91;
        399: twf_out = -118;
        400: twf_out = 128;
        401: twf_out = 126;
        402: twf_out = 118;
        403: twf_out = 106;
        404: twf_out = 91;
        405: twf_out = 71;
        406: twf_out = 49;
        407: twf_out = 25;
        408: twf_out = 128;
        409: twf_out = 106;
        410: twf_out = 49;
        411: twf_out = -25;
        412: twf_out = -91;
        413: twf_out = -126;
        414: twf_out = -118;
        415: twf_out = -71;
        416: twf_out = 128;
        417: twf_out = 127;
        418: twf_out = 126;
        419: twf_out = 122;
        420: twf_out = 118;
        421: twf_out = 113;
        422: twf_out = 106;
        423: twf_out = 99;
        424: twf_out = 128;
        425: twf_out = 113;
        426: twf_out = 71;
        427: twf_out = 13;
        428: twf_out = -49;
        429: twf_out = -99;
        430: twf_out = -126;
        431: twf_out = -122;
        432: twf_out = 128;
        433: twf_out = 122;
        434: twf_out = 106;
        435: twf_out = 81;
        436: twf_out = 49;
        437: twf_out = 13;
        438: twf_out = -25;
        439: twf_out = -60;
        440: twf_out = 128;
        441: twf_out = 99;
        442: twf_out = 25;
        443: twf_out = -60;
        444: twf_out = -118;
        445: twf_out = -122;
        446: twf_out = -71;
        447: twf_out = 13;
        448: twf_out = 128;
        449: twf_out = 128;
        450: twf_out = 128;
        451: twf_out = 128;
        452: twf_out = 128;
        453: twf_out = 128;
        454: twf_out = 128;
        455: twf_out = 128;
        456: twf_out = 128;
        457: twf_out = 118;
        458: twf_out = 91;
        459: twf_out = 49;
        460: twf_out = 0;
        461: twf_out = -49;
        462: twf_out = -91;
        463: twf_out = -118;
        464: twf_out = 128;
        465: twf_out = 126;
        466: twf_out = 118;
        467: twf_out = 106;
        468: twf_out = 91;
        469: twf_out = 71;
        470: twf_out = 49;
        471: twf_out = 25;
        472: twf_out = 128;
        473: twf_out = 106;
        474: twf_out = 49;
        475: twf_out = -25;
        476: twf_out = -91;
        477: twf_out = -126;
        478: twf_out = -118;
        479: twf_out = -71;
        480: twf_out = 128;
        481: twf_out = 127;
        482: twf_out = 126;
        483: twf_out = 122;
        484: twf_out = 118;
        485: twf_out = 113;
        486: twf_out = 106;
        487: twf_out = 99;
        488: twf_out = 128;
        489: twf_out = 113;
        490: twf_out = 71;
        491: twf_out = 13;
        492: twf_out = -49;
        493: twf_out = -99;
        494: twf_out = -126;
        495: twf_out = -122;
        496: twf_out = 128;
        497: twf_out = 122;
        498: twf_out = 106;
        499: twf_out = 81;
        500: twf_out = 49;
        501: twf_out = 13;
        502: twf_out = -25;
        503: twf_out = -60;
        504: twf_out = 128;
        505: twf_out = 99;
        506: twf_out = 25;
        507: twf_out = -60;
        508: twf_out = -118;
        509: twf_out = -122;
        510: twf_out = -71;
        511: twf_out = 13;
        default: twf_out = 0;
    endcase
end

endmodule

`timescale 1ns/1ps

module step02_twf #(
    parameter INDEX_WIDTH = 512,
    parameter BIT_WIDTH = 9 //2.7format
) (
    input [$clog2(INDEX_WIDTH)-1:0] index,
    output signed [BIT_WIDTH-1:0] twf_out
);

wire signed [BIT_WIDTH-1:0] twf_02_out [0:INDEX_WIDTH-1];

assign twf_out = twf_02_out[index];

assign twf_02_out[0] = 128;
assign twf_02_out[1] = 128;
assign twf_02_out[2] = 128;
assign twf_02_out[3] = 128;
assign twf_02_out[4] = 128;
assign twf_02_out[5] = 128;
assign twf_02_out[6] = 128;
assign twf_02_out[7] = 128;
assign twf_02_out[8] = 128;
assign twf_02_out[9] = 128;
assign twf_02_out[10] = 128;
assign twf_02_out[11] = 128;
assign twf_02_out[12] = 128;
assign twf_02_out[13] = 128;
assign twf_02_out[14] = 128;
assign twf_02_out[15] = 128;
assign twf_02_out[16] = 128;
assign twf_02_out[17] = 128;
assign twf_02_out[18] = 128;
assign twf_02_out[19] = 128;
assign twf_02_out[20] = 128;
assign twf_02_out[21] = 128;
assign twf_02_out[22] = 128;
assign twf_02_out[23] = 128;
assign twf_02_out[24] = 128;
assign twf_02_out[25] = 128;
assign twf_02_out[26] = 128;
assign twf_02_out[27] = 128;
assign twf_02_out[28] = 128;
assign twf_02_out[29] = 128;
assign twf_02_out[30] = 128;
assign twf_02_out[31] = 128;
assign twf_02_out[32] = 128;
assign twf_02_out[33] = 128;
assign twf_02_out[34] = 128;
assign twf_02_out[35] = 128;
assign twf_02_out[36] = 128;
assign twf_02_out[37] = 128;
assign twf_02_out[38] = 128;
assign twf_02_out[39] = 128;
assign twf_02_out[40] = 128;
assign twf_02_out[41] = 128;
assign twf_02_out[42] = 128;
assign twf_02_out[43] = 128;
assign twf_02_out[44] = 128;
assign twf_02_out[45] = 128;
assign twf_02_out[46] = 128;
assign twf_02_out[47] = 128;
assign twf_02_out[48] = 128;
assign twf_02_out[49] = 128;
assign twf_02_out[50] = 128;
assign twf_02_out[51] = 128;
assign twf_02_out[52] = 128;
assign twf_02_out[53] = 128;
assign twf_02_out[54] = 128;
assign twf_02_out[55] = 128;
assign twf_02_out[56] = 128;
assign twf_02_out[57] = 128;
assign twf_02_out[58] = 128;
assign twf_02_out[59] = 128;
assign twf_02_out[60] = 128;
assign twf_02_out[61] = 128;
assign twf_02_out[62] = 128;
assign twf_02_out[63] = 128;
assign twf_02_out[64] = 128;
assign twf_02_out[65] = 128;
assign twf_02_out[66] = 127;
assign twf_02_out[67] = 127;
assign twf_02_out[68] = 126;
assign twf_02_out[69] = 124;
assign twf_02_out[70] = 122;
assign twf_02_out[71] = 121;
assign twf_02_out[72] = 118;
assign twf_02_out[73] = 116;
assign twf_02_out[74] = 113;
assign twf_02_out[75] = 110;
assign twf_02_out[76] = 106;
assign twf_02_out[77] = 103;
assign twf_02_out[78] = 99;
assign twf_02_out[79] = 95;
assign twf_02_out[80] = 91;
assign twf_02_out[81] = 86;
assign twf_02_out[82] = 81;
assign twf_02_out[83] = 76;
assign twf_02_out[84] = 71;
assign twf_02_out[85] = 66;
assign twf_02_out[86] = 60;
assign twf_02_out[87] = 55;
assign twf_02_out[88] = 49;
assign twf_02_out[89] = 43;
assign twf_02_out[90] = 37;
assign twf_02_out[91] = 31;
assign twf_02_out[92] = 25;
assign twf_02_out[93] = 19;
assign twf_02_out[94] = 13;
assign twf_02_out[95] = 6;
assign twf_02_out[96] = 0;
assign twf_02_out[97] = -6;
assign twf_02_out[98] = -13;
assign twf_02_out[99] = -19;
assign twf_02_out[100] = -25;
assign twf_02_out[101] = -31;
assign twf_02_out[102] = -37;
assign twf_02_out[103] = -43;
assign twf_02_out[104] = -49;
assign twf_02_out[105] = -55;
assign twf_02_out[106] = -60;
assign twf_02_out[107] = -66;
assign twf_02_out[108] = -71;
assign twf_02_out[109] = -76;
assign twf_02_out[110] = -81;
assign twf_02_out[111] = -86;
assign twf_02_out[112] = -91;
assign twf_02_out[113] = -95;
assign twf_02_out[114] = -99;
assign twf_02_out[115] = -103;
assign twf_02_out[116] = -106;
assign twf_02_out[117] = -110;
assign twf_02_out[118] = -113;
assign twf_02_out[119] = -116;
assign twf_02_out[120] = -118;
assign twf_02_out[121] = -121;
assign twf_02_out[122] = -122;
assign twf_02_out[123] = -124;
assign twf_02_out[124] = -126;
assign twf_02_out[125] = -127;
assign twf_02_out[126] = -127;
assign twf_02_out[127] = -128;
assign twf_02_out[128] = 128;
assign twf_02_out[129] = 128;
assign twf_02_out[130] = 128;
assign twf_02_out[131] = 128;
assign twf_02_out[132] = 127;
assign twf_02_out[133] = 127;
assign twf_02_out[134] = 127;
assign twf_02_out[135] = 126;
assign twf_02_out[136] = 126;
assign twf_02_out[137] = 125;
assign twf_02_out[138] = 124;
assign twf_02_out[139] = 123;
assign twf_02_out[140] = 122;
assign twf_02_out[141] = 122;
assign twf_02_out[142] = 121;
assign twf_02_out[143] = 119;
assign twf_02_out[144] = 118;
assign twf_02_out[145] = 117;
assign twf_02_out[146] = 116;
assign twf_02_out[147] = 114;
assign twf_02_out[148] = 113;
assign twf_02_out[149] = 111;
assign twf_02_out[150] = 110;
assign twf_02_out[151] = 108;
assign twf_02_out[152] = 106;
assign twf_02_out[153] = 105;
assign twf_02_out[154] = 103;
assign twf_02_out[155] = 101;
assign twf_02_out[156] = 99;
assign twf_02_out[157] = 97;
assign twf_02_out[158] = 95;
assign twf_02_out[159] = 93;
assign twf_02_out[160] = 91;
assign twf_02_out[161] = 88;
assign twf_02_out[162] = 86;
assign twf_02_out[163] = 84;
assign twf_02_out[164] = 81;
assign twf_02_out[165] = 79;
assign twf_02_out[166] = 76;
assign twf_02_out[167] = 74;
assign twf_02_out[168] = 71;
assign twf_02_out[169] = 68;
assign twf_02_out[170] = 66;
assign twf_02_out[171] = 63;
assign twf_02_out[172] = 60;
assign twf_02_out[173] = 58;
assign twf_02_out[174] = 55;
assign twf_02_out[175] = 52;
assign twf_02_out[176] = 49;
assign twf_02_out[177] = 46;
assign twf_02_out[178] = 43;
assign twf_02_out[179] = 40;
assign twf_02_out[180] = 37;
assign twf_02_out[181] = 34;
assign twf_02_out[182] = 31;
assign twf_02_out[183] = 28;
assign twf_02_out[184] = 25;
assign twf_02_out[185] = 22;
assign twf_02_out[186] = 19;
assign twf_02_out[187] = 16;
assign twf_02_out[188] = 13;
assign twf_02_out[189] = 9;
assign twf_02_out[190] = 6;
assign twf_02_out[191] = 3;
assign twf_02_out[192] = 128;
assign twf_02_out[193] = 128;
assign twf_02_out[194] = 127;
assign twf_02_out[195] = 125;
assign twf_02_out[196] = 122;
assign twf_02_out[197] = 119;
assign twf_02_out[198] = 116;
assign twf_02_out[199] = 111;
assign twf_02_out[200] = 106;
assign twf_02_out[201] = 101;
assign twf_02_out[202] = 95;
assign twf_02_out[203] = 88;
assign twf_02_out[204] = 81;
assign twf_02_out[205] = 74;
assign twf_02_out[206] = 66;
assign twf_02_out[207] = 58;
assign twf_02_out[208] = 49;
assign twf_02_out[209] = 40;
assign twf_02_out[210] = 31;
assign twf_02_out[211] = 22;
assign twf_02_out[212] = 13;
assign twf_02_out[213] = 3;
assign twf_02_out[214] = -6;
assign twf_02_out[215] = -16;
assign twf_02_out[216] = -25;
assign twf_02_out[217] = -34;
assign twf_02_out[218] = -43;
assign twf_02_out[219] = -52;
assign twf_02_out[220] = -60;
assign twf_02_out[221] = -68;
assign twf_02_out[222] = -76;
assign twf_02_out[223] = -84;
assign twf_02_out[224] = -91;
assign twf_02_out[225] = -97;
assign twf_02_out[226] = -103;
assign twf_02_out[227] = -108;
assign twf_02_out[228] = -113;
assign twf_02_out[229] = -117;
assign twf_02_out[230] = -121;
assign twf_02_out[231] = -123;
assign twf_02_out[232] = -126;
assign twf_02_out[233] = -127;
assign twf_02_out[234] = -128;
assign twf_02_out[235] = -128;
assign twf_02_out[236] = -127;
assign twf_02_out[237] = -126;
assign twf_02_out[238] = -124;
assign twf_02_out[239] = -122;
assign twf_02_out[240] = -118;
assign twf_02_out[241] = -114;
assign twf_02_out[242] = -110;
assign twf_02_out[243] = -105;
assign twf_02_out[244] = -99;
assign twf_02_out[245] = -93;
assign twf_02_out[246] = -86;
assign twf_02_out[247] = -79;
assign twf_02_out[248] = -71;
assign twf_02_out[249] = -63;
assign twf_02_out[250] = -55;
assign twf_02_out[251] = -46;
assign twf_02_out[252] = -37;
assign twf_02_out[253] = -28;
assign twf_02_out[254] = -19;
assign twf_02_out[255] = -9;
assign twf_02_out[256] = 128;
assign twf_02_out[257] = 128;
assign twf_02_out[258] = 128;
assign twf_02_out[259] = 128;
assign twf_02_out[260] = 128;
assign twf_02_out[261] = 128;
assign twf_02_out[262] = 128;
assign twf_02_out[263] = 128;
assign twf_02_out[264] = 127;
assign twf_02_out[265] = 127;
assign twf_02_out[266] = 127;
assign twf_02_out[267] = 127;
assign twf_02_out[268] = 127;
assign twf_02_out[269] = 126;
assign twf_02_out[270] = 126;
assign twf_02_out[271] = 126;
assign twf_02_out[272] = 126;
assign twf_02_out[273] = 125;
assign twf_02_out[274] = 125;
assign twf_02_out[275] = 125;
assign twf_02_out[276] = 124;
assign twf_02_out[277] = 124;
assign twf_02_out[278] = 123;
assign twf_02_out[279] = 123;
assign twf_02_out[280] = 122;
assign twf_02_out[281] = 122;
assign twf_02_out[282] = 122;
assign twf_02_out[283] = 121;
assign twf_02_out[284] = 121;
assign twf_02_out[285] = 120;
assign twf_02_out[286] = 119;
assign twf_02_out[287] = 119;
assign twf_02_out[288] = 118;
assign twf_02_out[289] = 118;
assign twf_02_out[290] = 117;
assign twf_02_out[291] = 116;
assign twf_02_out[292] = 116;
assign twf_02_out[293] = 115;
assign twf_02_out[294] = 114;
assign twf_02_out[295] = 114;
assign twf_02_out[296] = 113;
assign twf_02_out[297] = 112;
assign twf_02_out[298] = 111;
assign twf_02_out[299] = 111;
assign twf_02_out[300] = 110;
assign twf_02_out[301] = 109;
assign twf_02_out[302] = 108;
assign twf_02_out[303] = 107;
assign twf_02_out[304] = 106;
assign twf_02_out[305] = 106;
assign twf_02_out[306] = 105;
assign twf_02_out[307] = 104;
assign twf_02_out[308] = 103;
assign twf_02_out[309] = 102;
assign twf_02_out[310] = 101;
assign twf_02_out[311] = 100;
assign twf_02_out[312] = 99;
assign twf_02_out[313] = 98;
assign twf_02_out[314] = 97;
assign twf_02_out[315] = 96;
assign twf_02_out[316] = 95;
assign twf_02_out[317] = 94;
assign twf_02_out[318] = 93;
assign twf_02_out[319] = 92;
assign twf_02_out[320] = 128;
assign twf_02_out[321] = 128;
assign twf_02_out[322] = 127;
assign twf_02_out[323] = 126;
assign twf_02_out[324] = 124;
assign twf_02_out[325] = 122;
assign twf_02_out[326] = 119;
assign twf_02_out[327] = 116;
assign twf_02_out[328] = 113;
assign twf_02_out[329] = 109;
assign twf_02_out[330] = 105;
assign twf_02_out[331] = 100;
assign twf_02_out[332] = 95;
assign twf_02_out[333] = 89;
assign twf_02_out[334] = 84;
assign twf_02_out[335] = 78;
assign twf_02_out[336] = 71;
assign twf_02_out[337] = 64;
assign twf_02_out[338] = 58;
assign twf_02_out[339] = 50;
assign twf_02_out[340] = 43;
assign twf_02_out[341] = 36;
assign twf_02_out[342] = 28;
assign twf_02_out[343] = 20;
assign twf_02_out[344] = 13;
assign twf_02_out[345] = 5;
assign twf_02_out[346] = -3;
assign twf_02_out[347] = -11;
assign twf_02_out[348] = -19;
assign twf_02_out[349] = -27;
assign twf_02_out[350] = -34;
assign twf_02_out[351] = -42;
assign twf_02_out[352] = -49;
assign twf_02_out[353] = -56;
assign twf_02_out[354] = -63;
assign twf_02_out[355] = -70;
assign twf_02_out[356] = -76;
assign twf_02_out[357] = -82;
assign twf_02_out[358] = -88;
assign twf_02_out[359] = -94;
assign twf_02_out[360] = -99;
assign twf_02_out[361] = -104;
assign twf_02_out[362] = -108;
assign twf_02_out[363] = -112;
assign twf_02_out[364] = -116;
assign twf_02_out[365] = -119;
assign twf_02_out[366] = -122;
assign twf_02_out[367] = -124;
assign twf_02_out[368] = -126;
assign twf_02_out[369] = -127;
assign twf_02_out[370] = -128;
assign twf_02_out[371] = -128;
assign twf_02_out[372] = -128;
assign twf_02_out[373] = -127;
assign twf_02_out[374] = -126;
assign twf_02_out[375] = -125;
assign twf_02_out[376] = -122;
assign twf_02_out[377] = -120;
assign twf_02_out[378] = -117;
assign twf_02_out[379] = -114;
assign twf_02_out[380] = -110;
assign twf_02_out[381] = -106;
assign twf_02_out[382] = -101;
assign twf_02_out[383] = -96;
assign twf_02_out[384] = 128;
assign twf_02_out[385] = 128;
assign twf_02_out[386] = 128;
assign twf_02_out[387] = 127;
assign twf_02_out[388] = 127;
assign twf_02_out[389] = 126;
assign twf_02_out[390] = 125;
assign twf_02_out[391] = 124;
assign twf_02_out[392] = 122;
assign twf_02_out[393] = 121;
assign twf_02_out[394] = 119;
assign twf_02_out[395] = 118;
assign twf_02_out[396] = 116;
assign twf_02_out[397] = 114;
assign twf_02_out[398] = 111;
assign twf_02_out[399] = 109;
assign twf_02_out[400] = 106;
assign twf_02_out[401] = 104;
assign twf_02_out[402] = 101;
assign twf_02_out[403] = 98;
assign twf_02_out[404] = 95;
assign twf_02_out[405] = 92;
assign twf_02_out[406] = 88;
assign twf_02_out[407] = 85;
assign twf_02_out[408] = 81;
assign twf_02_out[409] = 78;
assign twf_02_out[410] = 74;
assign twf_02_out[411] = 70;
assign twf_02_out[412] = 66;
assign twf_02_out[413] = 62;
assign twf_02_out[414] = 58;
assign twf_02_out[415] = 53;
assign twf_02_out[416] = 49;
assign twf_02_out[417] = 45;
assign twf_02_out[418] = 40;
assign twf_02_out[419] = 36;
assign twf_02_out[420] = 31;
assign twf_02_out[421] = 27;
assign twf_02_out[422] = 22;
assign twf_02_out[423] = 17;
assign twf_02_out[424] = 13;
assign twf_02_out[425] = 8;
assign twf_02_out[426] = 3;
assign twf_02_out[427] = -2;
assign twf_02_out[428] = -6;
assign twf_02_out[429] = -11;
assign twf_02_out[430] = -16;
assign twf_02_out[431] = -20;
assign twf_02_out[432] = -25;
assign twf_02_out[433] = -30;
assign twf_02_out[434] = -34;
assign twf_02_out[435] = -39;
assign twf_02_out[436] = -43;
assign twf_02_out[437] = -48;
assign twf_02_out[438] = -52;
assign twf_02_out[439] = -56;
assign twf_02_out[440] = -60;
assign twf_02_out[441] = -64;
assign twf_02_out[442] = -68;
assign twf_02_out[443] = -72;
assign twf_02_out[444] = -76;
assign twf_02_out[445] = -80;
assign twf_02_out[446] = -84;
assign twf_02_out[447] = -87;
assign twf_02_out[448] = 128;
assign twf_02_out[449] = 128;
assign twf_02_out[450] = 126;
assign twf_02_out[451] = 124;
assign twf_02_out[452] = 121;
assign twf_02_out[453] = 116;
assign twf_02_out[454] = 111;
assign twf_02_out[455] = 106;
assign twf_02_out[456] = 99;
assign twf_02_out[457] = 92;
assign twf_02_out[458] = 84;
assign twf_02_out[459] = 75;
assign twf_02_out[460] = 66;
assign twf_02_out[461] = 56;
assign twf_02_out[462] = 46;
assign twf_02_out[463] = 36;
assign twf_02_out[464] = 25;
assign twf_02_out[465] = 14;
assign twf_02_out[466] = 3;
assign twf_02_out[467] = -8;
assign twf_02_out[468] = -19;
assign twf_02_out[469] = -30;
assign twf_02_out[470] = -40;
assign twf_02_out[471] = -50;
assign twf_02_out[472] = -60;
assign twf_02_out[473] = -70;
assign twf_02_out[474] = -79;
assign twf_02_out[475] = -87;
assign twf_02_out[476] = -95;
assign twf_02_out[477] = -102;
assign twf_02_out[478] = -108;
assign twf_02_out[479] = -114;
assign twf_02_out[480] = -118;
assign twf_02_out[481] = -122;
assign twf_02_out[482] = -125;
assign twf_02_out[483] = -127;
assign twf_02_out[484] = -128;
assign twf_02_out[485] = -128;
assign twf_02_out[486] = -127;
assign twf_02_out[487] = -125;
assign twf_02_out[488] = -122;
assign twf_02_out[489] = -119;
assign twf_02_out[490] = -114;
assign twf_02_out[491] = -109;
assign twf_02_out[492] = -103;
assign twf_02_out[493] = -96;
assign twf_02_out[494] = -88;
assign twf_02_out[495] = -80;
assign twf_02_out[496] = -71;
assign twf_02_out[497] = -62;
assign twf_02_out[498] = -52;
assign twf_02_out[499] = -42;
assign twf_02_out[500] = -31;
assign twf_02_out[501] = -20;
assign twf_02_out[502] = -9;
assign twf_02_out[503] = 2;
assign twf_02_out[504] = 13;
assign twf_02_out[505] = 23;
assign twf_02_out[506] = 34;
assign twf_02_out[507] = 45;
assign twf_02_out[508] = 55;
assign twf_02_out[509] = 64;
assign twf_02_out[510] = 74;
assign twf_02_out[511] = 82;

endmodule